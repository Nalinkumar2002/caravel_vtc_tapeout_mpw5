magic
tech sky130A
timestamp 1647751980
<< nwell >>
rect 19624 16012 20522 16014
rect 18761 15833 20630 16012
rect 17447 15228 17930 15630
rect 18759 15265 20630 15833
rect 17627 15227 17930 15228
rect 18767 15012 20630 15265
rect 19198 15011 20630 15012
rect 19422 15010 20630 15011
rect 17221 14009 18134 14382
rect 17453 14008 18043 14009
<< pwell >>
rect 17479 14788 17613 14986
rect 17291 14662 17613 14788
rect 17755 14788 17889 14985
rect 17291 14519 17425 14662
rect 17755 14661 18077 14788
rect 17943 14562 18077 14661
rect 17943 14519 18070 14562
rect 17284 14462 18070 14519
rect 18819 14438 18953 14946
rect 19249 14436 19383 14944
rect 19648 14717 19782 14943
rect 19716 14656 19782 14717
rect 19913 14656 20047 14945
rect 20183 14656 20317 14945
rect 20454 14717 20588 14943
rect 20454 14656 20502 14717
rect 19716 14599 20502 14656
rect 18963 14284 19219 14342
rect 17339 13420 17473 13846
rect 17887 13420 18021 13846
rect 17615 13035 17749 13333
rect 17564 12977 17820 13035
<< nmos >>
rect 17537 14873 17555 14973
rect 17813 14872 17831 14972
rect 17349 14575 17367 14775
rect 17537 14675 17555 14775
rect 17813 14674 17831 14774
rect 18001 14575 18019 14775
rect 18877 14733 18895 14933
rect 19307 14731 19325 14931
rect 19706 14730 19724 14930
rect 19971 14732 19989 14932
rect 20241 14732 20259 14932
rect 20512 14730 20530 14930
rect 18877 14451 18895 14651
rect 19307 14449 19325 14649
rect 17397 13433 17415 13833
rect 17945 13433 17963 13833
rect 17673 13120 17691 13320
<< pmos >>
rect 17537 15254 17555 15454
rect 17812 15253 17830 15453
rect 18875 15089 18893 15289
rect 19305 15087 19323 15287
rect 19706 15044 19724 15844
rect 19971 15046 19989 15846
rect 20241 15046 20259 15846
rect 20512 15044 20530 15844
rect 17397 14036 17415 14236
rect 17946 14034 17964 14234
<< ndiff >>
rect 17492 14957 17537 14973
rect 17492 14939 17501 14957
rect 17519 14939 17537 14957
rect 17492 14907 17537 14939
rect 17492 14889 17501 14907
rect 17519 14889 17537 14907
rect 17492 14873 17537 14889
rect 17555 14956 17600 14973
rect 17555 14938 17573 14956
rect 17591 14938 17600 14956
rect 17555 14907 17600 14938
rect 17555 14889 17573 14907
rect 17591 14889 17600 14907
rect 17555 14873 17600 14889
rect 17768 14956 17813 14972
rect 17768 14938 17777 14956
rect 17795 14938 17813 14956
rect 17768 14906 17813 14938
rect 17768 14888 17777 14906
rect 17795 14888 17813 14906
rect 17768 14872 17813 14888
rect 17831 14955 17876 14972
rect 17831 14937 17849 14955
rect 17867 14937 17876 14955
rect 17831 14906 17876 14937
rect 17831 14888 17849 14906
rect 17867 14888 17876 14906
rect 17831 14872 17876 14888
rect 18832 14923 18877 14933
rect 18832 14905 18841 14923
rect 18859 14905 18877 14923
rect 18832 14885 18877 14905
rect 18832 14867 18841 14885
rect 18859 14867 18877 14885
rect 18832 14847 18877 14867
rect 18832 14829 18841 14847
rect 18859 14829 18877 14847
rect 17304 14765 17349 14775
rect 17304 14747 17313 14765
rect 17331 14747 17349 14765
rect 17304 14727 17349 14747
rect 17304 14709 17313 14727
rect 17331 14709 17349 14727
rect 17304 14689 17349 14709
rect 17304 14671 17313 14689
rect 17331 14671 17349 14689
rect 17304 14650 17349 14671
rect 17304 14632 17313 14650
rect 17331 14632 17349 14650
rect 17304 14609 17349 14632
rect 17304 14591 17313 14609
rect 17331 14591 17349 14609
rect 17304 14575 17349 14591
rect 17367 14765 17412 14775
rect 17367 14747 17385 14765
rect 17403 14747 17412 14765
rect 17367 14727 17412 14747
rect 17367 14709 17385 14727
rect 17403 14709 17412 14727
rect 17367 14689 17412 14709
rect 17367 14671 17385 14689
rect 17403 14671 17412 14689
rect 17492 14759 17537 14775
rect 17492 14741 17501 14759
rect 17519 14741 17537 14759
rect 17492 14709 17537 14741
rect 17492 14691 17501 14709
rect 17519 14691 17537 14709
rect 17492 14675 17537 14691
rect 17555 14758 17600 14775
rect 18832 14808 18877 14829
rect 18832 14790 18841 14808
rect 18859 14790 18877 14808
rect 17555 14740 17573 14758
rect 17591 14740 17600 14758
rect 17555 14709 17600 14740
rect 17555 14691 17573 14709
rect 17591 14691 17600 14709
rect 17555 14675 17600 14691
rect 17768 14758 17813 14774
rect 17768 14740 17777 14758
rect 17795 14740 17813 14758
rect 17768 14708 17813 14740
rect 17768 14690 17777 14708
rect 17795 14690 17813 14708
rect 17367 14650 17412 14671
rect 17768 14674 17813 14690
rect 17831 14757 17876 14774
rect 17831 14739 17849 14757
rect 17867 14739 17876 14757
rect 17831 14708 17876 14739
rect 17831 14690 17849 14708
rect 17867 14690 17876 14708
rect 17831 14674 17876 14690
rect 17956 14765 18001 14775
rect 17956 14747 17965 14765
rect 17983 14747 18001 14765
rect 17956 14727 18001 14747
rect 17956 14709 17965 14727
rect 17983 14709 18001 14727
rect 17956 14689 18001 14709
rect 17956 14671 17965 14689
rect 17983 14671 18001 14689
rect 17367 14632 17385 14650
rect 17403 14632 17412 14650
rect 17367 14609 17412 14632
rect 17367 14591 17385 14609
rect 17403 14591 17412 14609
rect 17367 14575 17412 14591
rect 17956 14650 18001 14671
rect 17956 14632 17965 14650
rect 17983 14632 18001 14650
rect 17956 14609 18001 14632
rect 17956 14591 17965 14609
rect 17983 14591 18001 14609
rect 17956 14575 18001 14591
rect 18019 14765 18064 14775
rect 18019 14747 18037 14765
rect 18055 14747 18064 14765
rect 18019 14727 18064 14747
rect 18832 14767 18877 14790
rect 18832 14749 18841 14767
rect 18859 14749 18877 14767
rect 18832 14733 18877 14749
rect 18895 14923 18940 14933
rect 18895 14905 18913 14923
rect 18931 14905 18940 14923
rect 18895 14885 18940 14905
rect 18895 14867 18913 14885
rect 18931 14867 18940 14885
rect 18895 14847 18940 14867
rect 18895 14829 18913 14847
rect 18931 14829 18940 14847
rect 18895 14808 18940 14829
rect 18895 14790 18913 14808
rect 18931 14790 18940 14808
rect 18895 14767 18940 14790
rect 18895 14749 18913 14767
rect 18931 14749 18940 14767
rect 18895 14733 18940 14749
rect 19262 14921 19307 14931
rect 19262 14903 19271 14921
rect 19289 14903 19307 14921
rect 19262 14883 19307 14903
rect 19262 14865 19271 14883
rect 19289 14865 19307 14883
rect 19262 14845 19307 14865
rect 19262 14827 19271 14845
rect 19289 14827 19307 14845
rect 19262 14806 19307 14827
rect 19262 14788 19271 14806
rect 19289 14788 19307 14806
rect 19262 14765 19307 14788
rect 19262 14747 19271 14765
rect 19289 14747 19307 14765
rect 18019 14709 18037 14727
rect 18055 14709 18064 14727
rect 19262 14731 19307 14747
rect 19325 14921 19370 14931
rect 19325 14903 19343 14921
rect 19361 14903 19370 14921
rect 19325 14883 19370 14903
rect 19325 14865 19343 14883
rect 19361 14865 19370 14883
rect 19325 14845 19370 14865
rect 19325 14827 19343 14845
rect 19361 14827 19370 14845
rect 19325 14806 19370 14827
rect 19325 14788 19343 14806
rect 19361 14788 19370 14806
rect 19325 14765 19370 14788
rect 19325 14747 19343 14765
rect 19361 14747 19370 14765
rect 19325 14731 19370 14747
rect 19661 14920 19706 14930
rect 19661 14902 19670 14920
rect 19688 14902 19706 14920
rect 19661 14882 19706 14902
rect 19661 14864 19670 14882
rect 19688 14864 19706 14882
rect 19661 14844 19706 14864
rect 19661 14826 19670 14844
rect 19688 14826 19706 14844
rect 19661 14805 19706 14826
rect 19661 14787 19670 14805
rect 19688 14787 19706 14805
rect 19661 14764 19706 14787
rect 19661 14746 19670 14764
rect 19688 14746 19706 14764
rect 19661 14730 19706 14746
rect 19724 14920 19769 14930
rect 19724 14902 19742 14920
rect 19760 14902 19769 14920
rect 19724 14882 19769 14902
rect 19724 14864 19742 14882
rect 19760 14864 19769 14882
rect 19724 14844 19769 14864
rect 19724 14826 19742 14844
rect 19760 14826 19769 14844
rect 19724 14805 19769 14826
rect 19724 14787 19742 14805
rect 19760 14787 19769 14805
rect 19724 14764 19769 14787
rect 19724 14746 19742 14764
rect 19760 14746 19769 14764
rect 19724 14730 19769 14746
rect 19926 14922 19971 14932
rect 19926 14904 19935 14922
rect 19953 14904 19971 14922
rect 19926 14884 19971 14904
rect 19926 14866 19935 14884
rect 19953 14866 19971 14884
rect 19926 14846 19971 14866
rect 19926 14828 19935 14846
rect 19953 14828 19971 14846
rect 19926 14807 19971 14828
rect 19926 14789 19935 14807
rect 19953 14789 19971 14807
rect 19926 14766 19971 14789
rect 19926 14748 19935 14766
rect 19953 14748 19971 14766
rect 19926 14732 19971 14748
rect 19989 14922 20034 14932
rect 19989 14904 20007 14922
rect 20025 14904 20034 14922
rect 19989 14884 20034 14904
rect 19989 14866 20007 14884
rect 20025 14866 20034 14884
rect 19989 14846 20034 14866
rect 19989 14828 20007 14846
rect 20025 14828 20034 14846
rect 19989 14807 20034 14828
rect 19989 14789 20007 14807
rect 20025 14789 20034 14807
rect 19989 14766 20034 14789
rect 19989 14748 20007 14766
rect 20025 14748 20034 14766
rect 19989 14732 20034 14748
rect 20196 14922 20241 14932
rect 20196 14904 20205 14922
rect 20223 14904 20241 14922
rect 20196 14884 20241 14904
rect 20196 14866 20205 14884
rect 20223 14866 20241 14884
rect 20196 14846 20241 14866
rect 20196 14828 20205 14846
rect 20223 14828 20241 14846
rect 20196 14807 20241 14828
rect 20196 14789 20205 14807
rect 20223 14789 20241 14807
rect 20196 14766 20241 14789
rect 20196 14748 20205 14766
rect 20223 14748 20241 14766
rect 20196 14732 20241 14748
rect 20259 14922 20304 14932
rect 20259 14904 20277 14922
rect 20295 14904 20304 14922
rect 20259 14884 20304 14904
rect 20259 14866 20277 14884
rect 20295 14866 20304 14884
rect 20259 14846 20304 14866
rect 20259 14828 20277 14846
rect 20295 14828 20304 14846
rect 20259 14807 20304 14828
rect 20259 14789 20277 14807
rect 20295 14789 20304 14807
rect 20259 14766 20304 14789
rect 20259 14748 20277 14766
rect 20295 14748 20304 14766
rect 20259 14732 20304 14748
rect 20467 14920 20512 14930
rect 20467 14902 20476 14920
rect 20494 14902 20512 14920
rect 20467 14882 20512 14902
rect 20467 14864 20476 14882
rect 20494 14864 20512 14882
rect 20467 14844 20512 14864
rect 20467 14826 20476 14844
rect 20494 14826 20512 14844
rect 20467 14805 20512 14826
rect 20467 14787 20476 14805
rect 20494 14787 20512 14805
rect 20467 14764 20512 14787
rect 20467 14746 20476 14764
rect 20494 14746 20512 14764
rect 20467 14730 20512 14746
rect 20530 14920 20575 14930
rect 20530 14902 20548 14920
rect 20566 14902 20575 14920
rect 20530 14882 20575 14902
rect 20530 14864 20548 14882
rect 20566 14864 20575 14882
rect 20530 14844 20575 14864
rect 20530 14826 20548 14844
rect 20566 14826 20575 14844
rect 20530 14805 20575 14826
rect 20530 14787 20548 14805
rect 20566 14787 20575 14805
rect 20530 14764 20575 14787
rect 20530 14746 20548 14764
rect 20566 14746 20575 14764
rect 20530 14730 20575 14746
rect 18019 14689 18064 14709
rect 18019 14671 18037 14689
rect 18055 14671 18064 14689
rect 18019 14650 18064 14671
rect 18019 14632 18037 14650
rect 18055 14632 18064 14650
rect 18019 14609 18064 14632
rect 18019 14591 18037 14609
rect 18055 14591 18064 14609
rect 18019 14575 18064 14591
rect 18832 14635 18877 14651
rect 18832 14617 18841 14635
rect 18859 14617 18877 14635
rect 18832 14594 18877 14617
rect 18832 14576 18841 14594
rect 18859 14576 18877 14594
rect 18832 14555 18877 14576
rect 18832 14537 18841 14555
rect 18859 14537 18877 14555
rect 18832 14517 18877 14537
rect 18832 14499 18841 14517
rect 18859 14499 18877 14517
rect 18832 14479 18877 14499
rect 18832 14461 18841 14479
rect 18859 14461 18877 14479
rect 18832 14451 18877 14461
rect 18895 14635 18940 14651
rect 18895 14617 18913 14635
rect 18931 14617 18940 14635
rect 18895 14594 18940 14617
rect 18895 14576 18913 14594
rect 18931 14576 18940 14594
rect 18895 14555 18940 14576
rect 18895 14537 18913 14555
rect 18931 14537 18940 14555
rect 18895 14517 18940 14537
rect 18895 14499 18913 14517
rect 18931 14499 18940 14517
rect 18895 14479 18940 14499
rect 18895 14461 18913 14479
rect 18931 14461 18940 14479
rect 18895 14451 18940 14461
rect 19262 14633 19307 14649
rect 19262 14615 19271 14633
rect 19289 14615 19307 14633
rect 19262 14592 19307 14615
rect 19262 14574 19271 14592
rect 19289 14574 19307 14592
rect 19262 14553 19307 14574
rect 19262 14535 19271 14553
rect 19289 14535 19307 14553
rect 19262 14515 19307 14535
rect 19262 14497 19271 14515
rect 19289 14497 19307 14515
rect 19262 14477 19307 14497
rect 19262 14459 19271 14477
rect 19289 14459 19307 14477
rect 19262 14449 19307 14459
rect 19325 14633 19370 14649
rect 19325 14615 19343 14633
rect 19361 14615 19370 14633
rect 19325 14592 19370 14615
rect 19325 14574 19343 14592
rect 19361 14574 19370 14592
rect 19325 14553 19370 14574
rect 19325 14535 19343 14553
rect 19361 14535 19370 14553
rect 19325 14515 19370 14535
rect 19325 14497 19343 14515
rect 19361 14497 19370 14515
rect 19325 14477 19370 14497
rect 19325 14459 19343 14477
rect 19361 14459 19370 14477
rect 19325 14449 19370 14459
rect 17352 13823 17397 13833
rect 17352 13805 17361 13823
rect 17379 13805 17397 13823
rect 17352 13785 17397 13805
rect 17352 13767 17361 13785
rect 17379 13767 17397 13785
rect 17352 13747 17397 13767
rect 17352 13729 17361 13747
rect 17379 13729 17397 13747
rect 17352 13708 17397 13729
rect 17352 13690 17361 13708
rect 17379 13690 17397 13708
rect 17352 13664 17397 13690
rect 17352 13646 17361 13664
rect 17379 13646 17397 13664
rect 17352 13626 17397 13646
rect 17352 13608 17361 13626
rect 17379 13608 17397 13626
rect 17352 13585 17397 13608
rect 17352 13567 17361 13585
rect 17379 13567 17397 13585
rect 17352 13547 17397 13567
rect 17352 13529 17361 13547
rect 17379 13529 17397 13547
rect 17352 13508 17397 13529
rect 17352 13490 17361 13508
rect 17379 13490 17397 13508
rect 17352 13467 17397 13490
rect 17352 13449 17361 13467
rect 17379 13449 17397 13467
rect 17352 13433 17397 13449
rect 17415 13823 17460 13833
rect 17415 13805 17433 13823
rect 17451 13805 17460 13823
rect 17415 13785 17460 13805
rect 17415 13767 17433 13785
rect 17451 13767 17460 13785
rect 17415 13747 17460 13767
rect 17415 13729 17433 13747
rect 17451 13729 17460 13747
rect 17415 13708 17460 13729
rect 17415 13690 17433 13708
rect 17451 13690 17460 13708
rect 17415 13664 17460 13690
rect 17415 13646 17433 13664
rect 17451 13646 17460 13664
rect 17415 13626 17460 13646
rect 17415 13608 17433 13626
rect 17451 13608 17460 13626
rect 17415 13585 17460 13608
rect 17415 13567 17433 13585
rect 17451 13567 17460 13585
rect 17415 13547 17460 13567
rect 17415 13529 17433 13547
rect 17451 13529 17460 13547
rect 17415 13508 17460 13529
rect 17415 13490 17433 13508
rect 17451 13490 17460 13508
rect 17415 13467 17460 13490
rect 17415 13449 17433 13467
rect 17451 13449 17460 13467
rect 17415 13433 17460 13449
rect 17900 13823 17945 13833
rect 17900 13805 17909 13823
rect 17927 13805 17945 13823
rect 17900 13785 17945 13805
rect 17900 13767 17909 13785
rect 17927 13767 17945 13785
rect 17900 13747 17945 13767
rect 17900 13729 17909 13747
rect 17927 13729 17945 13747
rect 17900 13708 17945 13729
rect 17900 13690 17909 13708
rect 17927 13690 17945 13708
rect 17900 13664 17945 13690
rect 17900 13646 17909 13664
rect 17927 13646 17945 13664
rect 17900 13626 17945 13646
rect 17900 13608 17909 13626
rect 17927 13608 17945 13626
rect 17900 13585 17945 13608
rect 17900 13567 17909 13585
rect 17927 13567 17945 13585
rect 17900 13547 17945 13567
rect 17900 13529 17909 13547
rect 17927 13529 17945 13547
rect 17900 13508 17945 13529
rect 17900 13490 17909 13508
rect 17927 13490 17945 13508
rect 17900 13467 17945 13490
rect 17900 13449 17909 13467
rect 17927 13449 17945 13467
rect 17900 13433 17945 13449
rect 17963 13823 18008 13833
rect 17963 13805 17981 13823
rect 17999 13805 18008 13823
rect 17963 13785 18008 13805
rect 17963 13767 17981 13785
rect 17999 13767 18008 13785
rect 17963 13747 18008 13767
rect 17963 13729 17981 13747
rect 17999 13729 18008 13747
rect 17963 13708 18008 13729
rect 17963 13690 17981 13708
rect 17999 13690 18008 13708
rect 17963 13664 18008 13690
rect 17963 13646 17981 13664
rect 17999 13646 18008 13664
rect 17963 13626 18008 13646
rect 17963 13608 17981 13626
rect 17999 13608 18008 13626
rect 17963 13585 18008 13608
rect 17963 13567 17981 13585
rect 17999 13567 18008 13585
rect 17963 13547 18008 13567
rect 17963 13529 17981 13547
rect 17999 13529 18008 13547
rect 17963 13508 18008 13529
rect 17963 13490 17981 13508
rect 17999 13490 18008 13508
rect 17963 13467 18008 13490
rect 17963 13449 17981 13467
rect 17999 13449 18008 13467
rect 17963 13433 18008 13449
rect 17628 13310 17673 13320
rect 17628 13292 17637 13310
rect 17655 13292 17673 13310
rect 17628 13272 17673 13292
rect 17628 13254 17637 13272
rect 17655 13254 17673 13272
rect 17628 13234 17673 13254
rect 17628 13216 17637 13234
rect 17655 13216 17673 13234
rect 17628 13195 17673 13216
rect 17628 13177 17637 13195
rect 17655 13177 17673 13195
rect 17628 13154 17673 13177
rect 17628 13136 17637 13154
rect 17655 13136 17673 13154
rect 17628 13120 17673 13136
rect 17691 13310 17736 13320
rect 17691 13292 17709 13310
rect 17727 13292 17736 13310
rect 17691 13272 17736 13292
rect 17691 13254 17709 13272
rect 17727 13254 17736 13272
rect 17691 13234 17736 13254
rect 17691 13216 17709 13234
rect 17727 13216 17736 13234
rect 17691 13195 17736 13216
rect 17691 13177 17709 13195
rect 17727 13177 17736 13195
rect 17691 13154 17736 13177
rect 17691 13136 17709 13154
rect 17727 13136 17736 13154
rect 17691 13120 17736 13136
<< pdiff >>
rect 19661 15828 19706 15844
rect 19661 15810 19670 15828
rect 19688 15810 19706 15828
rect 19661 15787 19706 15810
rect 19661 15769 19670 15787
rect 19688 15769 19706 15787
rect 19661 15748 19706 15769
rect 19661 15730 19670 15748
rect 19688 15730 19706 15748
rect 19661 15710 19706 15730
rect 19661 15692 19670 15710
rect 19688 15692 19706 15710
rect 19661 15672 19706 15692
rect 19661 15654 19670 15672
rect 19688 15654 19706 15672
rect 19661 15628 19706 15654
rect 19661 15610 19670 15628
rect 19688 15610 19706 15628
rect 19661 15587 19706 15610
rect 19661 15569 19670 15587
rect 19688 15569 19706 15587
rect 19661 15548 19706 15569
rect 19661 15530 19670 15548
rect 19688 15530 19706 15548
rect 19661 15510 19706 15530
rect 19661 15492 19670 15510
rect 19688 15492 19706 15510
rect 19661 15472 19706 15492
rect 17492 15444 17537 15454
rect 17492 15426 17501 15444
rect 17519 15426 17537 15444
rect 17492 15406 17537 15426
rect 17492 15388 17501 15406
rect 17519 15388 17537 15406
rect 17492 15368 17537 15388
rect 17492 15350 17501 15368
rect 17519 15350 17537 15368
rect 17492 15329 17537 15350
rect 17492 15311 17501 15329
rect 17519 15311 17537 15329
rect 17492 15288 17537 15311
rect 17492 15270 17501 15288
rect 17519 15270 17537 15288
rect 17492 15254 17537 15270
rect 17555 15444 17600 15454
rect 19661 15454 19670 15472
rect 19688 15454 19706 15472
rect 17555 15426 17573 15444
rect 17591 15426 17600 15444
rect 17555 15406 17600 15426
rect 17555 15388 17573 15406
rect 17591 15388 17600 15406
rect 17555 15368 17600 15388
rect 17555 15350 17573 15368
rect 17591 15350 17600 15368
rect 17555 15329 17600 15350
rect 17555 15311 17573 15329
rect 17591 15311 17600 15329
rect 17555 15288 17600 15311
rect 17555 15270 17573 15288
rect 17591 15270 17600 15288
rect 17555 15254 17600 15270
rect 17767 15443 17812 15453
rect 17767 15425 17776 15443
rect 17794 15425 17812 15443
rect 17767 15405 17812 15425
rect 17767 15387 17776 15405
rect 17794 15387 17812 15405
rect 17767 15367 17812 15387
rect 17767 15349 17776 15367
rect 17794 15349 17812 15367
rect 17767 15328 17812 15349
rect 17767 15310 17776 15328
rect 17794 15310 17812 15328
rect 17767 15287 17812 15310
rect 17767 15269 17776 15287
rect 17794 15269 17812 15287
rect 17767 15253 17812 15269
rect 17830 15443 17875 15453
rect 17830 15425 17848 15443
rect 17866 15425 17875 15443
rect 17830 15405 17875 15425
rect 17830 15387 17848 15405
rect 17866 15387 17875 15405
rect 19661 15428 19706 15454
rect 19661 15410 19670 15428
rect 19688 15410 19706 15428
rect 17830 15367 17875 15387
rect 19661 15387 19706 15410
rect 17830 15349 17848 15367
rect 17866 15349 17875 15367
rect 17830 15328 17875 15349
rect 17830 15310 17848 15328
rect 17866 15310 17875 15328
rect 17830 15287 17875 15310
rect 19661 15369 19670 15387
rect 19688 15369 19706 15387
rect 19661 15348 19706 15369
rect 19661 15330 19670 15348
rect 19688 15330 19706 15348
rect 19661 15310 19706 15330
rect 17830 15269 17848 15287
rect 17866 15269 17875 15287
rect 17830 15253 17875 15269
rect 18830 15273 18875 15289
rect 18830 15255 18839 15273
rect 18857 15255 18875 15273
rect 18830 15232 18875 15255
rect 18830 15214 18839 15232
rect 18857 15214 18875 15232
rect 18830 15193 18875 15214
rect 18830 15175 18839 15193
rect 18857 15175 18875 15193
rect 18830 15155 18875 15175
rect 18830 15137 18839 15155
rect 18857 15137 18875 15155
rect 18830 15117 18875 15137
rect 18830 15099 18839 15117
rect 18857 15099 18875 15117
rect 18830 15089 18875 15099
rect 18893 15273 18938 15289
rect 19661 15292 19670 15310
rect 19688 15292 19706 15310
rect 18893 15255 18911 15273
rect 18929 15255 18938 15273
rect 18893 15232 18938 15255
rect 18893 15214 18911 15232
rect 18929 15214 18938 15232
rect 18893 15193 18938 15214
rect 18893 15175 18911 15193
rect 18929 15175 18938 15193
rect 18893 15155 18938 15175
rect 18893 15137 18911 15155
rect 18929 15137 18938 15155
rect 18893 15117 18938 15137
rect 18893 15099 18911 15117
rect 18929 15099 18938 15117
rect 18893 15089 18938 15099
rect 19260 15271 19305 15287
rect 19260 15253 19269 15271
rect 19287 15253 19305 15271
rect 19260 15230 19305 15253
rect 19260 15212 19269 15230
rect 19287 15212 19305 15230
rect 19260 15191 19305 15212
rect 19260 15173 19269 15191
rect 19287 15173 19305 15191
rect 19260 15153 19305 15173
rect 19260 15135 19269 15153
rect 19287 15135 19305 15153
rect 19260 15115 19305 15135
rect 19260 15097 19269 15115
rect 19287 15097 19305 15115
rect 19260 15087 19305 15097
rect 19323 15271 19368 15287
rect 19323 15253 19341 15271
rect 19359 15253 19368 15271
rect 19323 15230 19368 15253
rect 19323 15212 19341 15230
rect 19359 15212 19368 15230
rect 19323 15191 19368 15212
rect 19323 15173 19341 15191
rect 19359 15173 19368 15191
rect 19323 15153 19368 15173
rect 19323 15135 19341 15153
rect 19359 15135 19368 15153
rect 19323 15115 19368 15135
rect 19323 15097 19341 15115
rect 19359 15097 19368 15115
rect 19323 15087 19368 15097
rect 19661 15272 19706 15292
rect 19661 15254 19670 15272
rect 19688 15254 19706 15272
rect 19661 15228 19706 15254
rect 19661 15210 19670 15228
rect 19688 15210 19706 15228
rect 19661 15187 19706 15210
rect 19661 15169 19670 15187
rect 19688 15169 19706 15187
rect 19661 15148 19706 15169
rect 19661 15130 19670 15148
rect 19688 15130 19706 15148
rect 19661 15110 19706 15130
rect 19661 15092 19670 15110
rect 19688 15092 19706 15110
rect 19661 15072 19706 15092
rect 19661 15054 19670 15072
rect 19688 15054 19706 15072
rect 19661 15044 19706 15054
rect 19724 15828 19769 15844
rect 19724 15810 19742 15828
rect 19760 15810 19769 15828
rect 19724 15787 19769 15810
rect 19724 15769 19742 15787
rect 19760 15769 19769 15787
rect 19724 15748 19769 15769
rect 19724 15730 19742 15748
rect 19760 15730 19769 15748
rect 19724 15710 19769 15730
rect 19724 15692 19742 15710
rect 19760 15692 19769 15710
rect 19724 15672 19769 15692
rect 19724 15654 19742 15672
rect 19760 15654 19769 15672
rect 19724 15628 19769 15654
rect 19724 15610 19742 15628
rect 19760 15610 19769 15628
rect 19724 15587 19769 15610
rect 19724 15569 19742 15587
rect 19760 15569 19769 15587
rect 19724 15548 19769 15569
rect 19724 15530 19742 15548
rect 19760 15530 19769 15548
rect 19724 15510 19769 15530
rect 19724 15492 19742 15510
rect 19760 15492 19769 15510
rect 19724 15472 19769 15492
rect 19724 15454 19742 15472
rect 19760 15454 19769 15472
rect 19724 15428 19769 15454
rect 19724 15410 19742 15428
rect 19760 15410 19769 15428
rect 19724 15387 19769 15410
rect 19724 15369 19742 15387
rect 19760 15369 19769 15387
rect 19724 15348 19769 15369
rect 19724 15330 19742 15348
rect 19760 15330 19769 15348
rect 19724 15310 19769 15330
rect 19724 15292 19742 15310
rect 19760 15292 19769 15310
rect 19724 15272 19769 15292
rect 19724 15254 19742 15272
rect 19760 15254 19769 15272
rect 19724 15228 19769 15254
rect 19724 15210 19742 15228
rect 19760 15210 19769 15228
rect 19724 15187 19769 15210
rect 19724 15169 19742 15187
rect 19760 15169 19769 15187
rect 19724 15148 19769 15169
rect 19724 15130 19742 15148
rect 19760 15130 19769 15148
rect 19724 15110 19769 15130
rect 19724 15092 19742 15110
rect 19760 15092 19769 15110
rect 19724 15072 19769 15092
rect 19724 15054 19742 15072
rect 19760 15054 19769 15072
rect 19724 15044 19769 15054
rect 19926 15830 19971 15846
rect 19926 15812 19935 15830
rect 19953 15812 19971 15830
rect 19926 15789 19971 15812
rect 19926 15771 19935 15789
rect 19953 15771 19971 15789
rect 19926 15750 19971 15771
rect 19926 15732 19935 15750
rect 19953 15732 19971 15750
rect 19926 15712 19971 15732
rect 19926 15694 19935 15712
rect 19953 15694 19971 15712
rect 19926 15674 19971 15694
rect 19926 15656 19935 15674
rect 19953 15656 19971 15674
rect 19926 15630 19971 15656
rect 19926 15612 19935 15630
rect 19953 15612 19971 15630
rect 19926 15589 19971 15612
rect 19926 15571 19935 15589
rect 19953 15571 19971 15589
rect 19926 15550 19971 15571
rect 19926 15532 19935 15550
rect 19953 15532 19971 15550
rect 19926 15512 19971 15532
rect 19926 15494 19935 15512
rect 19953 15494 19971 15512
rect 19926 15474 19971 15494
rect 19926 15456 19935 15474
rect 19953 15456 19971 15474
rect 19926 15430 19971 15456
rect 19926 15412 19935 15430
rect 19953 15412 19971 15430
rect 19926 15389 19971 15412
rect 19926 15371 19935 15389
rect 19953 15371 19971 15389
rect 19926 15350 19971 15371
rect 19926 15332 19935 15350
rect 19953 15332 19971 15350
rect 19926 15312 19971 15332
rect 19926 15294 19935 15312
rect 19953 15294 19971 15312
rect 19926 15274 19971 15294
rect 19926 15256 19935 15274
rect 19953 15256 19971 15274
rect 19926 15230 19971 15256
rect 19926 15212 19935 15230
rect 19953 15212 19971 15230
rect 19926 15189 19971 15212
rect 19926 15171 19935 15189
rect 19953 15171 19971 15189
rect 19926 15150 19971 15171
rect 19926 15132 19935 15150
rect 19953 15132 19971 15150
rect 19926 15112 19971 15132
rect 19926 15094 19935 15112
rect 19953 15094 19971 15112
rect 19926 15074 19971 15094
rect 19926 15056 19935 15074
rect 19953 15056 19971 15074
rect 19926 15046 19971 15056
rect 19989 15830 20034 15846
rect 19989 15812 20007 15830
rect 20025 15812 20034 15830
rect 19989 15789 20034 15812
rect 19989 15771 20007 15789
rect 20025 15771 20034 15789
rect 19989 15750 20034 15771
rect 19989 15732 20007 15750
rect 20025 15732 20034 15750
rect 19989 15712 20034 15732
rect 19989 15694 20007 15712
rect 20025 15694 20034 15712
rect 19989 15674 20034 15694
rect 19989 15656 20007 15674
rect 20025 15656 20034 15674
rect 19989 15630 20034 15656
rect 19989 15612 20007 15630
rect 20025 15612 20034 15630
rect 19989 15589 20034 15612
rect 19989 15571 20007 15589
rect 20025 15571 20034 15589
rect 19989 15550 20034 15571
rect 19989 15532 20007 15550
rect 20025 15532 20034 15550
rect 19989 15512 20034 15532
rect 19989 15494 20007 15512
rect 20025 15494 20034 15512
rect 19989 15474 20034 15494
rect 19989 15456 20007 15474
rect 20025 15456 20034 15474
rect 19989 15430 20034 15456
rect 19989 15412 20007 15430
rect 20025 15412 20034 15430
rect 19989 15389 20034 15412
rect 19989 15371 20007 15389
rect 20025 15371 20034 15389
rect 19989 15350 20034 15371
rect 19989 15332 20007 15350
rect 20025 15332 20034 15350
rect 19989 15312 20034 15332
rect 19989 15294 20007 15312
rect 20025 15294 20034 15312
rect 19989 15274 20034 15294
rect 19989 15256 20007 15274
rect 20025 15256 20034 15274
rect 19989 15230 20034 15256
rect 19989 15212 20007 15230
rect 20025 15212 20034 15230
rect 19989 15189 20034 15212
rect 19989 15171 20007 15189
rect 20025 15171 20034 15189
rect 19989 15150 20034 15171
rect 19989 15132 20007 15150
rect 20025 15132 20034 15150
rect 19989 15112 20034 15132
rect 19989 15094 20007 15112
rect 20025 15094 20034 15112
rect 19989 15074 20034 15094
rect 19989 15056 20007 15074
rect 20025 15056 20034 15074
rect 19989 15046 20034 15056
rect 20196 15830 20241 15846
rect 20196 15812 20205 15830
rect 20223 15812 20241 15830
rect 20196 15789 20241 15812
rect 20196 15771 20205 15789
rect 20223 15771 20241 15789
rect 20196 15750 20241 15771
rect 20196 15732 20205 15750
rect 20223 15732 20241 15750
rect 20196 15712 20241 15732
rect 20196 15694 20205 15712
rect 20223 15694 20241 15712
rect 20196 15674 20241 15694
rect 20196 15656 20205 15674
rect 20223 15656 20241 15674
rect 20196 15630 20241 15656
rect 20196 15612 20205 15630
rect 20223 15612 20241 15630
rect 20196 15589 20241 15612
rect 20196 15571 20205 15589
rect 20223 15571 20241 15589
rect 20196 15550 20241 15571
rect 20196 15532 20205 15550
rect 20223 15532 20241 15550
rect 20196 15512 20241 15532
rect 20196 15494 20205 15512
rect 20223 15494 20241 15512
rect 20196 15474 20241 15494
rect 20196 15456 20205 15474
rect 20223 15456 20241 15474
rect 20196 15430 20241 15456
rect 20196 15412 20205 15430
rect 20223 15412 20241 15430
rect 20196 15389 20241 15412
rect 20196 15371 20205 15389
rect 20223 15371 20241 15389
rect 20196 15350 20241 15371
rect 20196 15332 20205 15350
rect 20223 15332 20241 15350
rect 20196 15312 20241 15332
rect 20196 15294 20205 15312
rect 20223 15294 20241 15312
rect 20196 15274 20241 15294
rect 20196 15256 20205 15274
rect 20223 15256 20241 15274
rect 20196 15230 20241 15256
rect 20196 15212 20205 15230
rect 20223 15212 20241 15230
rect 20196 15189 20241 15212
rect 20196 15171 20205 15189
rect 20223 15171 20241 15189
rect 20196 15150 20241 15171
rect 20196 15132 20205 15150
rect 20223 15132 20241 15150
rect 20196 15112 20241 15132
rect 20196 15094 20205 15112
rect 20223 15094 20241 15112
rect 20196 15074 20241 15094
rect 20196 15056 20205 15074
rect 20223 15056 20241 15074
rect 20196 15046 20241 15056
rect 20259 15830 20304 15846
rect 20259 15812 20277 15830
rect 20295 15812 20304 15830
rect 20259 15789 20304 15812
rect 20259 15771 20277 15789
rect 20295 15771 20304 15789
rect 20259 15750 20304 15771
rect 20259 15732 20277 15750
rect 20295 15732 20304 15750
rect 20259 15712 20304 15732
rect 20259 15694 20277 15712
rect 20295 15694 20304 15712
rect 20259 15674 20304 15694
rect 20259 15656 20277 15674
rect 20295 15656 20304 15674
rect 20259 15630 20304 15656
rect 20259 15612 20277 15630
rect 20295 15612 20304 15630
rect 20259 15589 20304 15612
rect 20259 15571 20277 15589
rect 20295 15571 20304 15589
rect 20259 15550 20304 15571
rect 20259 15532 20277 15550
rect 20295 15532 20304 15550
rect 20259 15512 20304 15532
rect 20259 15494 20277 15512
rect 20295 15494 20304 15512
rect 20259 15474 20304 15494
rect 20259 15456 20277 15474
rect 20295 15456 20304 15474
rect 20259 15430 20304 15456
rect 20259 15412 20277 15430
rect 20295 15412 20304 15430
rect 20259 15389 20304 15412
rect 20259 15371 20277 15389
rect 20295 15371 20304 15389
rect 20259 15350 20304 15371
rect 20259 15332 20277 15350
rect 20295 15332 20304 15350
rect 20259 15312 20304 15332
rect 20259 15294 20277 15312
rect 20295 15294 20304 15312
rect 20259 15274 20304 15294
rect 20259 15256 20277 15274
rect 20295 15256 20304 15274
rect 20259 15230 20304 15256
rect 20259 15212 20277 15230
rect 20295 15212 20304 15230
rect 20259 15189 20304 15212
rect 20259 15171 20277 15189
rect 20295 15171 20304 15189
rect 20259 15150 20304 15171
rect 20259 15132 20277 15150
rect 20295 15132 20304 15150
rect 20259 15112 20304 15132
rect 20259 15094 20277 15112
rect 20295 15094 20304 15112
rect 20259 15074 20304 15094
rect 20259 15056 20277 15074
rect 20295 15056 20304 15074
rect 20259 15046 20304 15056
rect 20467 15828 20512 15844
rect 20467 15810 20476 15828
rect 20494 15810 20512 15828
rect 20467 15787 20512 15810
rect 20467 15769 20476 15787
rect 20494 15769 20512 15787
rect 20467 15748 20512 15769
rect 20467 15730 20476 15748
rect 20494 15730 20512 15748
rect 20467 15710 20512 15730
rect 20467 15692 20476 15710
rect 20494 15692 20512 15710
rect 20467 15672 20512 15692
rect 20467 15654 20476 15672
rect 20494 15654 20512 15672
rect 20467 15628 20512 15654
rect 20467 15610 20476 15628
rect 20494 15610 20512 15628
rect 20467 15587 20512 15610
rect 20467 15569 20476 15587
rect 20494 15569 20512 15587
rect 20467 15548 20512 15569
rect 20467 15530 20476 15548
rect 20494 15530 20512 15548
rect 20467 15510 20512 15530
rect 20467 15492 20476 15510
rect 20494 15492 20512 15510
rect 20467 15472 20512 15492
rect 20467 15454 20476 15472
rect 20494 15454 20512 15472
rect 20467 15428 20512 15454
rect 20467 15410 20476 15428
rect 20494 15410 20512 15428
rect 20467 15387 20512 15410
rect 20467 15369 20476 15387
rect 20494 15369 20512 15387
rect 20467 15348 20512 15369
rect 20467 15330 20476 15348
rect 20494 15330 20512 15348
rect 20467 15310 20512 15330
rect 20467 15292 20476 15310
rect 20494 15292 20512 15310
rect 20467 15272 20512 15292
rect 20467 15254 20476 15272
rect 20494 15254 20512 15272
rect 20467 15228 20512 15254
rect 20467 15210 20476 15228
rect 20494 15210 20512 15228
rect 20467 15187 20512 15210
rect 20467 15169 20476 15187
rect 20494 15169 20512 15187
rect 20467 15148 20512 15169
rect 20467 15130 20476 15148
rect 20494 15130 20512 15148
rect 20467 15110 20512 15130
rect 20467 15092 20476 15110
rect 20494 15092 20512 15110
rect 20467 15072 20512 15092
rect 20467 15054 20476 15072
rect 20494 15054 20512 15072
rect 20467 15044 20512 15054
rect 20530 15828 20575 15844
rect 20530 15810 20548 15828
rect 20566 15810 20575 15828
rect 20530 15787 20575 15810
rect 20530 15769 20548 15787
rect 20566 15769 20575 15787
rect 20530 15748 20575 15769
rect 20530 15730 20548 15748
rect 20566 15730 20575 15748
rect 20530 15710 20575 15730
rect 20530 15692 20548 15710
rect 20566 15692 20575 15710
rect 20530 15672 20575 15692
rect 20530 15654 20548 15672
rect 20566 15654 20575 15672
rect 20530 15628 20575 15654
rect 20530 15610 20548 15628
rect 20566 15610 20575 15628
rect 20530 15587 20575 15610
rect 20530 15569 20548 15587
rect 20566 15569 20575 15587
rect 20530 15548 20575 15569
rect 20530 15530 20548 15548
rect 20566 15530 20575 15548
rect 20530 15510 20575 15530
rect 20530 15492 20548 15510
rect 20566 15492 20575 15510
rect 20530 15472 20575 15492
rect 20530 15454 20548 15472
rect 20566 15454 20575 15472
rect 20530 15428 20575 15454
rect 20530 15410 20548 15428
rect 20566 15410 20575 15428
rect 20530 15387 20575 15410
rect 20530 15369 20548 15387
rect 20566 15369 20575 15387
rect 20530 15348 20575 15369
rect 20530 15330 20548 15348
rect 20566 15330 20575 15348
rect 20530 15310 20575 15330
rect 20530 15292 20548 15310
rect 20566 15292 20575 15310
rect 20530 15272 20575 15292
rect 20530 15254 20548 15272
rect 20566 15254 20575 15272
rect 20530 15228 20575 15254
rect 20530 15210 20548 15228
rect 20566 15210 20575 15228
rect 20530 15187 20575 15210
rect 20530 15169 20548 15187
rect 20566 15169 20575 15187
rect 20530 15148 20575 15169
rect 20530 15130 20548 15148
rect 20566 15130 20575 15148
rect 20530 15110 20575 15130
rect 20530 15092 20548 15110
rect 20566 15092 20575 15110
rect 20530 15072 20575 15092
rect 20530 15054 20548 15072
rect 20566 15054 20575 15072
rect 20530 15044 20575 15054
rect 17352 14226 17397 14236
rect 17352 14208 17361 14226
rect 17379 14208 17397 14226
rect 17352 14188 17397 14208
rect 17352 14170 17361 14188
rect 17379 14170 17397 14188
rect 17352 14150 17397 14170
rect 17352 14132 17361 14150
rect 17379 14132 17397 14150
rect 17352 14111 17397 14132
rect 17352 14093 17361 14111
rect 17379 14093 17397 14111
rect 17352 14070 17397 14093
rect 17352 14052 17361 14070
rect 17379 14052 17397 14070
rect 17352 14036 17397 14052
rect 17415 14226 17460 14236
rect 17415 14208 17433 14226
rect 17451 14208 17460 14226
rect 17415 14188 17460 14208
rect 17415 14170 17433 14188
rect 17451 14170 17460 14188
rect 17415 14150 17460 14170
rect 17415 14132 17433 14150
rect 17451 14132 17460 14150
rect 17415 14111 17460 14132
rect 17415 14093 17433 14111
rect 17451 14093 17460 14111
rect 17415 14070 17460 14093
rect 17415 14052 17433 14070
rect 17451 14052 17460 14070
rect 17415 14036 17460 14052
rect 17901 14224 17946 14234
rect 17901 14206 17910 14224
rect 17928 14206 17946 14224
rect 17901 14186 17946 14206
rect 17901 14168 17910 14186
rect 17928 14168 17946 14186
rect 17901 14148 17946 14168
rect 17901 14130 17910 14148
rect 17928 14130 17946 14148
rect 17901 14109 17946 14130
rect 17901 14091 17910 14109
rect 17928 14091 17946 14109
rect 17901 14068 17946 14091
rect 17901 14050 17910 14068
rect 17928 14050 17946 14068
rect 17901 14034 17946 14050
rect 17964 14224 18009 14234
rect 17964 14206 17982 14224
rect 18000 14206 18009 14224
rect 17964 14186 18009 14206
rect 17964 14168 17982 14186
rect 18000 14168 18009 14186
rect 17964 14148 18009 14168
rect 17964 14130 17982 14148
rect 18000 14130 18009 14148
rect 17964 14109 18009 14130
rect 17964 14091 17982 14109
rect 18000 14091 18009 14109
rect 17964 14068 18009 14091
rect 17964 14050 17982 14068
rect 18000 14050 18009 14068
rect 17964 14034 18009 14050
<< ndiffc >>
rect 17501 14939 17519 14957
rect 17501 14889 17519 14907
rect 17573 14938 17591 14956
rect 17573 14889 17591 14907
rect 17777 14938 17795 14956
rect 17777 14888 17795 14906
rect 17849 14937 17867 14955
rect 17849 14888 17867 14906
rect 18841 14905 18859 14923
rect 18841 14867 18859 14885
rect 18841 14829 18859 14847
rect 17313 14747 17331 14765
rect 17313 14709 17331 14727
rect 17313 14671 17331 14689
rect 17313 14632 17331 14650
rect 17313 14591 17331 14609
rect 17385 14747 17403 14765
rect 17385 14709 17403 14727
rect 17385 14671 17403 14689
rect 17501 14741 17519 14759
rect 17501 14691 17519 14709
rect 18841 14790 18859 14808
rect 17573 14740 17591 14758
rect 17573 14691 17591 14709
rect 17777 14740 17795 14758
rect 17777 14690 17795 14708
rect 17849 14739 17867 14757
rect 17849 14690 17867 14708
rect 17965 14747 17983 14765
rect 17965 14709 17983 14727
rect 17965 14671 17983 14689
rect 17385 14632 17403 14650
rect 17385 14591 17403 14609
rect 17965 14632 17983 14650
rect 17965 14591 17983 14609
rect 18037 14747 18055 14765
rect 18841 14749 18859 14767
rect 18913 14905 18931 14923
rect 18913 14867 18931 14885
rect 18913 14829 18931 14847
rect 18913 14790 18931 14808
rect 18913 14749 18931 14767
rect 19271 14903 19289 14921
rect 19271 14865 19289 14883
rect 19271 14827 19289 14845
rect 19271 14788 19289 14806
rect 19271 14747 19289 14765
rect 18037 14709 18055 14727
rect 19343 14903 19361 14921
rect 19343 14865 19361 14883
rect 19343 14827 19361 14845
rect 19343 14788 19361 14806
rect 19343 14747 19361 14765
rect 19670 14902 19688 14920
rect 19670 14864 19688 14882
rect 19670 14826 19688 14844
rect 19670 14787 19688 14805
rect 19670 14746 19688 14764
rect 19742 14902 19760 14920
rect 19742 14864 19760 14882
rect 19742 14826 19760 14844
rect 19742 14787 19760 14805
rect 19742 14746 19760 14764
rect 19935 14904 19953 14922
rect 19935 14866 19953 14884
rect 19935 14828 19953 14846
rect 19935 14789 19953 14807
rect 19935 14748 19953 14766
rect 20007 14904 20025 14922
rect 20007 14866 20025 14884
rect 20007 14828 20025 14846
rect 20007 14789 20025 14807
rect 20007 14748 20025 14766
rect 20205 14904 20223 14922
rect 20205 14866 20223 14884
rect 20205 14828 20223 14846
rect 20205 14789 20223 14807
rect 20205 14748 20223 14766
rect 20277 14904 20295 14922
rect 20277 14866 20295 14884
rect 20277 14828 20295 14846
rect 20277 14789 20295 14807
rect 20277 14748 20295 14766
rect 20476 14902 20494 14920
rect 20476 14864 20494 14882
rect 20476 14826 20494 14844
rect 20476 14787 20494 14805
rect 20476 14746 20494 14764
rect 20548 14902 20566 14920
rect 20548 14864 20566 14882
rect 20548 14826 20566 14844
rect 20548 14787 20566 14805
rect 20548 14746 20566 14764
rect 18037 14671 18055 14689
rect 18037 14632 18055 14650
rect 18037 14591 18055 14609
rect 18841 14617 18859 14635
rect 18841 14576 18859 14594
rect 18841 14537 18859 14555
rect 18841 14499 18859 14517
rect 18841 14461 18859 14479
rect 18913 14617 18931 14635
rect 18913 14576 18931 14594
rect 18913 14537 18931 14555
rect 18913 14499 18931 14517
rect 18913 14461 18931 14479
rect 19271 14615 19289 14633
rect 19271 14574 19289 14592
rect 19271 14535 19289 14553
rect 19271 14497 19289 14515
rect 19271 14459 19289 14477
rect 19343 14615 19361 14633
rect 19343 14574 19361 14592
rect 19343 14535 19361 14553
rect 19343 14497 19361 14515
rect 19343 14459 19361 14477
rect 17361 13805 17379 13823
rect 17361 13767 17379 13785
rect 17361 13729 17379 13747
rect 17361 13690 17379 13708
rect 17361 13646 17379 13664
rect 17361 13608 17379 13626
rect 17361 13567 17379 13585
rect 17361 13529 17379 13547
rect 17361 13490 17379 13508
rect 17361 13449 17379 13467
rect 17433 13805 17451 13823
rect 17433 13767 17451 13785
rect 17433 13729 17451 13747
rect 17433 13690 17451 13708
rect 17433 13646 17451 13664
rect 17433 13608 17451 13626
rect 17433 13567 17451 13585
rect 17433 13529 17451 13547
rect 17433 13490 17451 13508
rect 17433 13449 17451 13467
rect 17909 13805 17927 13823
rect 17909 13767 17927 13785
rect 17909 13729 17927 13747
rect 17909 13690 17927 13708
rect 17909 13646 17927 13664
rect 17909 13608 17927 13626
rect 17909 13567 17927 13585
rect 17909 13529 17927 13547
rect 17909 13490 17927 13508
rect 17909 13449 17927 13467
rect 17981 13805 17999 13823
rect 17981 13767 17999 13785
rect 17981 13729 17999 13747
rect 17981 13690 17999 13708
rect 17981 13646 17999 13664
rect 17981 13608 17999 13626
rect 17981 13567 17999 13585
rect 17981 13529 17999 13547
rect 17981 13490 17999 13508
rect 17981 13449 17999 13467
rect 17637 13292 17655 13310
rect 17637 13254 17655 13272
rect 17637 13216 17655 13234
rect 17637 13177 17655 13195
rect 17637 13136 17655 13154
rect 17709 13292 17727 13310
rect 17709 13254 17727 13272
rect 17709 13216 17727 13234
rect 17709 13177 17727 13195
rect 17709 13136 17727 13154
<< pdiffc >>
rect 19670 15810 19688 15828
rect 19670 15769 19688 15787
rect 19670 15730 19688 15748
rect 19670 15692 19688 15710
rect 19670 15654 19688 15672
rect 19670 15610 19688 15628
rect 19670 15569 19688 15587
rect 19670 15530 19688 15548
rect 19670 15492 19688 15510
rect 17501 15426 17519 15444
rect 17501 15388 17519 15406
rect 17501 15350 17519 15368
rect 17501 15311 17519 15329
rect 17501 15270 17519 15288
rect 19670 15454 19688 15472
rect 17573 15426 17591 15444
rect 17573 15388 17591 15406
rect 17573 15350 17591 15368
rect 17573 15311 17591 15329
rect 17573 15270 17591 15288
rect 17776 15425 17794 15443
rect 17776 15387 17794 15405
rect 17776 15349 17794 15367
rect 17776 15310 17794 15328
rect 17776 15269 17794 15287
rect 17848 15425 17866 15443
rect 17848 15387 17866 15405
rect 19670 15410 19688 15428
rect 17848 15349 17866 15367
rect 17848 15310 17866 15328
rect 19670 15369 19688 15387
rect 19670 15330 19688 15348
rect 17848 15269 17866 15287
rect 18839 15255 18857 15273
rect 18839 15214 18857 15232
rect 18839 15175 18857 15193
rect 18839 15137 18857 15155
rect 18839 15099 18857 15117
rect 19670 15292 19688 15310
rect 18911 15255 18929 15273
rect 18911 15214 18929 15232
rect 18911 15175 18929 15193
rect 18911 15137 18929 15155
rect 18911 15099 18929 15117
rect 19269 15253 19287 15271
rect 19269 15212 19287 15230
rect 19269 15173 19287 15191
rect 19269 15135 19287 15153
rect 19269 15097 19287 15115
rect 19341 15253 19359 15271
rect 19341 15212 19359 15230
rect 19341 15173 19359 15191
rect 19341 15135 19359 15153
rect 19341 15097 19359 15115
rect 19670 15254 19688 15272
rect 19670 15210 19688 15228
rect 19670 15169 19688 15187
rect 19670 15130 19688 15148
rect 19670 15092 19688 15110
rect 19670 15054 19688 15072
rect 19742 15810 19760 15828
rect 19742 15769 19760 15787
rect 19742 15730 19760 15748
rect 19742 15692 19760 15710
rect 19742 15654 19760 15672
rect 19742 15610 19760 15628
rect 19742 15569 19760 15587
rect 19742 15530 19760 15548
rect 19742 15492 19760 15510
rect 19742 15454 19760 15472
rect 19742 15410 19760 15428
rect 19742 15369 19760 15387
rect 19742 15330 19760 15348
rect 19742 15292 19760 15310
rect 19742 15254 19760 15272
rect 19742 15210 19760 15228
rect 19742 15169 19760 15187
rect 19742 15130 19760 15148
rect 19742 15092 19760 15110
rect 19742 15054 19760 15072
rect 19935 15812 19953 15830
rect 19935 15771 19953 15789
rect 19935 15732 19953 15750
rect 19935 15694 19953 15712
rect 19935 15656 19953 15674
rect 19935 15612 19953 15630
rect 19935 15571 19953 15589
rect 19935 15532 19953 15550
rect 19935 15494 19953 15512
rect 19935 15456 19953 15474
rect 19935 15412 19953 15430
rect 19935 15371 19953 15389
rect 19935 15332 19953 15350
rect 19935 15294 19953 15312
rect 19935 15256 19953 15274
rect 19935 15212 19953 15230
rect 19935 15171 19953 15189
rect 19935 15132 19953 15150
rect 19935 15094 19953 15112
rect 19935 15056 19953 15074
rect 20007 15812 20025 15830
rect 20007 15771 20025 15789
rect 20007 15732 20025 15750
rect 20007 15694 20025 15712
rect 20007 15656 20025 15674
rect 20007 15612 20025 15630
rect 20007 15571 20025 15589
rect 20007 15532 20025 15550
rect 20007 15494 20025 15512
rect 20007 15456 20025 15474
rect 20007 15412 20025 15430
rect 20007 15371 20025 15389
rect 20007 15332 20025 15350
rect 20007 15294 20025 15312
rect 20007 15256 20025 15274
rect 20007 15212 20025 15230
rect 20007 15171 20025 15189
rect 20007 15132 20025 15150
rect 20007 15094 20025 15112
rect 20007 15056 20025 15074
rect 20205 15812 20223 15830
rect 20205 15771 20223 15789
rect 20205 15732 20223 15750
rect 20205 15694 20223 15712
rect 20205 15656 20223 15674
rect 20205 15612 20223 15630
rect 20205 15571 20223 15589
rect 20205 15532 20223 15550
rect 20205 15494 20223 15512
rect 20205 15456 20223 15474
rect 20205 15412 20223 15430
rect 20205 15371 20223 15389
rect 20205 15332 20223 15350
rect 20205 15294 20223 15312
rect 20205 15256 20223 15274
rect 20205 15212 20223 15230
rect 20205 15171 20223 15189
rect 20205 15132 20223 15150
rect 20205 15094 20223 15112
rect 20205 15056 20223 15074
rect 20277 15812 20295 15830
rect 20277 15771 20295 15789
rect 20277 15732 20295 15750
rect 20277 15694 20295 15712
rect 20277 15656 20295 15674
rect 20277 15612 20295 15630
rect 20277 15571 20295 15589
rect 20277 15532 20295 15550
rect 20277 15494 20295 15512
rect 20277 15456 20295 15474
rect 20277 15412 20295 15430
rect 20277 15371 20295 15389
rect 20277 15332 20295 15350
rect 20277 15294 20295 15312
rect 20277 15256 20295 15274
rect 20277 15212 20295 15230
rect 20277 15171 20295 15189
rect 20277 15132 20295 15150
rect 20277 15094 20295 15112
rect 20277 15056 20295 15074
rect 20476 15810 20494 15828
rect 20476 15769 20494 15787
rect 20476 15730 20494 15748
rect 20476 15692 20494 15710
rect 20476 15654 20494 15672
rect 20476 15610 20494 15628
rect 20476 15569 20494 15587
rect 20476 15530 20494 15548
rect 20476 15492 20494 15510
rect 20476 15454 20494 15472
rect 20476 15410 20494 15428
rect 20476 15369 20494 15387
rect 20476 15330 20494 15348
rect 20476 15292 20494 15310
rect 20476 15254 20494 15272
rect 20476 15210 20494 15228
rect 20476 15169 20494 15187
rect 20476 15130 20494 15148
rect 20476 15092 20494 15110
rect 20476 15054 20494 15072
rect 20548 15810 20566 15828
rect 20548 15769 20566 15787
rect 20548 15730 20566 15748
rect 20548 15692 20566 15710
rect 20548 15654 20566 15672
rect 20548 15610 20566 15628
rect 20548 15569 20566 15587
rect 20548 15530 20566 15548
rect 20548 15492 20566 15510
rect 20548 15454 20566 15472
rect 20548 15410 20566 15428
rect 20548 15369 20566 15387
rect 20548 15330 20566 15348
rect 20548 15292 20566 15310
rect 20548 15254 20566 15272
rect 20548 15210 20566 15228
rect 20548 15169 20566 15187
rect 20548 15130 20566 15148
rect 20548 15092 20566 15110
rect 20548 15054 20566 15072
rect 17361 14208 17379 14226
rect 17361 14170 17379 14188
rect 17361 14132 17379 14150
rect 17361 14093 17379 14111
rect 17361 14052 17379 14070
rect 17433 14208 17451 14226
rect 17433 14170 17451 14188
rect 17433 14132 17451 14150
rect 17433 14093 17451 14111
rect 17433 14052 17451 14070
rect 17910 14206 17928 14224
rect 17910 14168 17928 14186
rect 17910 14130 17928 14148
rect 17910 14091 17928 14109
rect 17910 14050 17928 14068
rect 17982 14206 18000 14224
rect 17982 14168 18000 14186
rect 17982 14130 18000 14148
rect 17982 14091 18000 14109
rect 17982 14050 18000 14068
<< psubdiff >>
rect 17297 14500 18057 14506
rect 17297 14482 17366 14500
rect 17384 14482 17463 14500
rect 17481 14482 17553 14500
rect 17571 14482 17654 14500
rect 17672 14482 17751 14500
rect 17769 14482 17841 14500
rect 17859 14482 17926 14500
rect 17944 14482 18003 14500
rect 18021 14482 18057 14500
rect 17297 14475 18057 14482
rect 19729 14637 20489 14643
rect 19729 14619 19798 14637
rect 19816 14619 19895 14637
rect 19913 14619 19985 14637
rect 20003 14619 20086 14637
rect 20104 14619 20183 14637
rect 20201 14619 20273 14637
rect 20291 14619 20358 14637
rect 20376 14619 20435 14637
rect 20453 14619 20489 14637
rect 19729 14612 20489 14619
rect 18976 14323 19206 14329
rect 18976 14305 18988 14323
rect 19006 14305 19085 14323
rect 19103 14305 19175 14323
rect 19193 14305 19206 14323
rect 18976 14297 19206 14305
rect 17577 13016 17807 13022
rect 17577 12998 17589 13016
rect 17607 12998 17686 13016
rect 17704 12998 17776 13016
rect 17794 12998 17807 13016
rect 17577 12990 17807 12998
<< nsubdiff >>
rect 19653 15955 20368 15956
rect 19653 15950 20496 15955
rect 19653 15932 19715 15950
rect 19733 15949 20096 15950
rect 19733 15932 19936 15949
rect 19653 15931 19936 15932
rect 19954 15932 20096 15949
rect 20114 15932 20193 15950
rect 20211 15932 20405 15950
rect 20423 15932 20496 15950
rect 19954 15931 20496 15932
rect 19653 15925 20496 15931
rect 19874 15924 20032 15925
rect 20355 15924 20496 15925
rect 17468 15593 17909 15599
rect 17468 15575 17530 15593
rect 17548 15575 17637 15593
rect 17655 15575 17734 15593
rect 17752 15575 17824 15593
rect 17842 15575 17909 15593
rect 17468 15568 17909 15575
rect 18864 15396 19305 15402
rect 18864 15378 18926 15396
rect 18944 15378 19033 15396
rect 19051 15378 19130 15396
rect 19148 15378 19220 15396
rect 19238 15378 19305 15396
rect 18864 15371 19305 15378
rect 17261 14338 18115 14344
rect 17261 14320 17323 14338
rect 17341 14320 17430 14338
rect 17448 14320 17527 14338
rect 17545 14320 17617 14338
rect 17635 14320 17750 14338
rect 17768 14320 17857 14338
rect 17875 14320 17954 14338
rect 17972 14320 18044 14338
rect 18062 14320 18115 14338
rect 17261 14313 18115 14320
<< psubdiffcont >>
rect 17366 14482 17384 14500
rect 17463 14482 17481 14500
rect 17553 14482 17571 14500
rect 17654 14482 17672 14500
rect 17751 14482 17769 14500
rect 17841 14482 17859 14500
rect 17926 14482 17944 14500
rect 18003 14482 18021 14500
rect 19798 14619 19816 14637
rect 19895 14619 19913 14637
rect 19985 14619 20003 14637
rect 20086 14619 20104 14637
rect 20183 14619 20201 14637
rect 20273 14619 20291 14637
rect 20358 14619 20376 14637
rect 20435 14619 20453 14637
rect 18988 14305 19006 14323
rect 19085 14305 19103 14323
rect 19175 14305 19193 14323
rect 17589 12998 17607 13016
rect 17686 12998 17704 13016
rect 17776 12998 17794 13016
<< nsubdiffcont >>
rect 19715 15932 19733 15950
rect 19936 15931 19954 15949
rect 20096 15932 20114 15950
rect 20193 15932 20211 15950
rect 20405 15932 20423 15950
rect 17530 15575 17548 15593
rect 17637 15575 17655 15593
rect 17734 15575 17752 15593
rect 17824 15575 17842 15593
rect 18926 15378 18944 15396
rect 19033 15378 19051 15396
rect 19130 15378 19148 15396
rect 19220 15378 19238 15396
rect 17323 14320 17341 14338
rect 17430 14320 17448 14338
rect 17527 14320 17545 14338
rect 17617 14320 17635 14338
rect 17750 14320 17768 14338
rect 17857 14320 17875 14338
rect 17954 14320 17972 14338
rect 18044 14320 18062 14338
<< poly >>
rect 19706 15844 19724 15869
rect 19971 15846 19989 15871
rect 20241 15846 20259 15871
rect 17537 15454 17555 15467
rect 17812 15453 17830 15466
rect 17537 15221 17555 15254
rect 18875 15289 18893 15302
rect 17527 15211 17563 15221
rect 17812 15217 17830 15253
rect 17527 15193 17537 15211
rect 17554 15193 17563 15211
rect 17527 15184 17563 15193
rect 17797 15209 17849 15217
rect 17797 15191 17812 15209
rect 17830 15191 17849 15209
rect 17797 15182 17849 15191
rect 19305 15287 19323 15300
rect 18875 15074 18893 15089
rect 18841 15065 18893 15074
rect 19305 15072 19323 15087
rect 18841 15047 18849 15065
rect 18867 15047 18893 15065
rect 18841 15038 18893 15047
rect 19271 15063 19323 15072
rect 19271 15045 19279 15063
rect 19297 15045 19323 15063
rect 19271 15036 19323 15045
rect 20512 15844 20530 15869
rect 17529 15017 17563 15026
rect 17529 14999 17537 15017
rect 17555 14999 17563 15017
rect 17529 14990 17563 14999
rect 17805 15016 17839 15025
rect 17805 14998 17813 15016
rect 17831 14998 17839 15016
rect 19706 14998 19724 15044
rect 19971 15000 19989 15046
rect 20241 15000 20259 15046
rect 17537 14973 17555 14990
rect 17805 14989 17839 14998
rect 19672 14989 19724 14998
rect 17813 14972 17831 14989
rect 18843 14975 18895 14984
rect 17537 14860 17555 14873
rect 18843 14957 18851 14975
rect 18869 14957 18895 14975
rect 18843 14948 18895 14957
rect 18877 14933 18895 14948
rect 19273 14973 19325 14982
rect 19273 14955 19281 14973
rect 19299 14955 19325 14973
rect 19672 14971 19680 14989
rect 19698 14971 19724 14989
rect 19672 14962 19724 14971
rect 19937 14991 19989 15000
rect 19937 14973 19945 14991
rect 19963 14973 19989 14991
rect 19937 14964 19989 14973
rect 20207 14991 20259 15000
rect 20512 14998 20530 15044
rect 20207 14973 20215 14991
rect 20233 14973 20259 14991
rect 20207 14964 20259 14973
rect 19273 14946 19325 14955
rect 17813 14859 17831 14872
rect 17315 14817 17367 14826
rect 17315 14799 17323 14817
rect 17341 14799 17367 14817
rect 17315 14790 17367 14799
rect 17349 14775 17367 14790
rect 17537 14819 17590 14828
rect 17537 14801 17562 14819
rect 17580 14801 17590 14819
rect 17537 14792 17590 14801
rect 17779 14819 17831 14828
rect 17779 14801 17787 14819
rect 17805 14801 17831 14819
rect 17779 14792 17831 14801
rect 17537 14775 17555 14792
rect 17813 14774 17831 14792
rect 18001 14818 18053 14827
rect 18001 14800 18027 14818
rect 18045 14800 18053 14818
rect 18001 14791 18053 14800
rect 18001 14775 18019 14791
rect 17537 14662 17555 14675
rect 17813 14661 17831 14674
rect 19307 14931 19325 14946
rect 18877 14720 18895 14733
rect 19706 14930 19724 14962
rect 19971 14932 19989 14964
rect 20241 14932 20259 14964
rect 20478 14989 20530 14998
rect 20478 14971 20486 14989
rect 20504 14971 20530 14989
rect 20478 14962 20530 14971
rect 19307 14718 19325 14731
rect 20512 14930 20530 14962
rect 19706 14717 19724 14730
rect 19971 14719 19989 14732
rect 20241 14719 20259 14732
rect 20512 14717 20530 14730
rect 18877 14651 18895 14664
rect 17349 14562 17367 14575
rect 18001 14562 18019 14575
rect 19307 14649 19325 14662
rect 18877 14436 18895 14451
rect 18843 14427 18895 14436
rect 19307 14434 19325 14449
rect 18843 14409 18851 14427
rect 18869 14409 18895 14427
rect 18843 14400 18895 14409
rect 19273 14425 19325 14434
rect 19273 14407 19281 14425
rect 19299 14407 19325 14425
rect 19273 14398 19325 14407
rect 17397 14236 17415 14249
rect 17946 14234 17964 14247
rect 17397 14007 17415 14036
rect 17363 13998 17415 14007
rect 17363 13980 17371 13998
rect 17389 13980 17415 13998
rect 17363 13971 17415 13980
rect 17946 14003 17964 14034
rect 17946 13994 17998 14003
rect 17946 13976 17972 13994
rect 17990 13976 17998 13994
rect 17946 13967 17998 13976
rect 17363 13876 17415 13885
rect 17363 13858 17371 13876
rect 17389 13858 17415 13876
rect 17363 13849 17415 13858
rect 17397 13833 17415 13849
rect 17945 13876 17997 13885
rect 17945 13858 17971 13876
rect 17989 13858 17997 13876
rect 17945 13849 17997 13858
rect 17945 13833 17963 13849
rect 17397 13420 17415 13433
rect 17945 13420 17963 13433
rect 17673 13320 17691 13333
rect 17673 13098 17691 13120
rect 17639 13089 17691 13098
rect 17639 13071 17647 13089
rect 17665 13071 17691 13089
rect 17639 13062 17691 13071
<< polycont >>
rect 17537 15193 17554 15211
rect 17812 15191 17830 15209
rect 18849 15047 18867 15065
rect 19279 15045 19297 15063
rect 17537 14999 17555 15017
rect 17813 14998 17831 15016
rect 18851 14957 18869 14975
rect 19281 14955 19299 14973
rect 19680 14971 19698 14989
rect 19945 14973 19963 14991
rect 20215 14973 20233 14991
rect 17323 14799 17341 14817
rect 17562 14801 17580 14819
rect 17787 14801 17805 14819
rect 18027 14800 18045 14818
rect 20486 14971 20504 14989
rect 18851 14409 18869 14427
rect 19281 14407 19299 14425
rect 17371 13980 17389 13998
rect 17972 13976 17990 13994
rect 17371 13858 17389 13876
rect 17971 13858 17989 13876
rect 17647 13071 17665 13089
<< locali >>
rect 16223 17003 16312 17026
rect 16223 16985 16256 17003
rect 16273 16985 16312 17003
rect 16223 16964 16312 16985
rect 16256 13876 16274 16964
rect 22295 16151 22357 16184
rect 21811 16134 22316 16151
rect 22334 16134 22357 16151
rect 21811 16133 22357 16134
rect 19644 15956 19811 15957
rect 19644 15955 20368 15956
rect 19644 15952 20496 15955
rect 19431 15950 20496 15952
rect 19431 15932 19669 15950
rect 19687 15932 19715 15950
rect 19733 15932 19769 15950
rect 19787 15949 20096 15950
rect 19787 15932 19890 15949
rect 19431 15931 19890 15932
rect 19908 15931 19936 15949
rect 19954 15931 19990 15949
rect 20008 15932 20096 15949
rect 20114 15932 20147 15950
rect 20165 15932 20193 15950
rect 20211 15932 20361 15950
rect 20379 15932 20405 15950
rect 20423 15932 20448 15950
rect 20466 15932 20496 15950
rect 20008 15931 20496 15932
rect 19431 15925 20496 15931
rect 19431 15924 20032 15925
rect 17468 15598 17909 15599
rect 17161 15593 18702 15598
rect 17161 15575 17484 15593
rect 17502 15575 17530 15593
rect 17548 15575 17584 15593
rect 17602 15575 17637 15593
rect 17655 15575 17688 15593
rect 17706 15575 17734 15593
rect 17752 15575 17780 15593
rect 17798 15575 17824 15593
rect 17842 15575 17867 15593
rect 17885 15575 18702 15593
rect 17161 15568 18702 15575
rect 17161 15567 17520 15568
rect 17102 15020 17136 15029
rect 17102 15002 17110 15020
rect 17128 15002 17136 15020
rect 17102 14993 17136 15002
rect 17044 14815 17075 14834
rect 17044 14798 17051 14815
rect 17068 14798 17075 14815
rect 17044 14778 17075 14798
rect 17045 13949 17063 14778
rect 17161 14344 17192 15567
rect 17501 15452 17519 15567
rect 17493 15444 17527 15452
rect 17493 15426 17501 15444
rect 17519 15426 17527 15444
rect 17493 15406 17527 15426
rect 17493 15388 17501 15406
rect 17519 15388 17527 15406
rect 17493 15368 17527 15388
rect 17493 15350 17501 15368
rect 17519 15350 17527 15368
rect 17493 15329 17527 15350
rect 17493 15311 17501 15329
rect 17519 15311 17527 15329
rect 17493 15288 17527 15311
rect 17493 15270 17501 15288
rect 17519 15270 17527 15288
rect 17493 15255 17527 15270
rect 17565 15444 17599 15453
rect 17848 15452 17866 15568
rect 17981 15566 18702 15568
rect 17565 15426 17573 15444
rect 17591 15426 17599 15444
rect 17565 15406 17599 15426
rect 17565 15388 17573 15406
rect 17591 15388 17599 15406
rect 17565 15368 17599 15388
rect 17565 15350 17573 15368
rect 17591 15350 17599 15368
rect 17565 15329 17599 15350
rect 17565 15311 17573 15329
rect 17591 15311 17599 15329
rect 17565 15288 17599 15311
rect 17768 15443 17802 15451
rect 17768 15425 17776 15443
rect 17794 15425 17802 15443
rect 17768 15405 17802 15425
rect 17768 15387 17776 15405
rect 17794 15387 17802 15405
rect 17768 15367 17802 15387
rect 17768 15349 17776 15367
rect 17794 15349 17802 15367
rect 17768 15328 17802 15349
rect 17768 15310 17776 15328
rect 17794 15310 17802 15328
rect 17565 15270 17573 15288
rect 17591 15270 17636 15288
rect 17768 15287 17802 15310
rect 17565 15255 17599 15270
rect 17527 15211 17563 15221
rect 17527 15193 17537 15211
rect 17554 15193 17563 15211
rect 17527 15184 17563 15193
rect 17370 15095 17422 15103
rect 17370 15077 17385 15095
rect 17403 15077 17422 15095
rect 17370 15068 17422 15077
rect 17618 15074 17636 15270
rect 17732 15269 17776 15287
rect 17794 15269 17802 15287
rect 17385 14834 17403 15068
rect 17607 15064 17643 15074
rect 17607 15046 17617 15064
rect 17634 15046 17643 15064
rect 17607 15037 17643 15046
rect 17529 15017 17563 15026
rect 17529 14999 17537 15017
rect 17555 14999 17563 15017
rect 17529 14990 17563 14999
rect 17493 14957 17527 14973
rect 17493 14939 17501 14957
rect 17519 14939 17527 14957
rect 17493 14907 17527 14939
rect 17493 14889 17501 14907
rect 17519 14889 17527 14907
rect 17493 14874 17527 14889
rect 17565 14956 17599 14973
rect 17618 14956 17636 15037
rect 17732 14956 17750 15269
rect 17768 15254 17802 15269
rect 17840 15443 17874 15452
rect 17840 15425 17848 15443
rect 17866 15425 17874 15443
rect 17840 15405 17874 15425
rect 17840 15387 17848 15405
rect 17866 15387 17874 15405
rect 17840 15367 17874 15387
rect 17840 15349 17848 15367
rect 17866 15349 17874 15367
rect 17840 15328 17874 15349
rect 17840 15310 17848 15328
rect 17866 15310 17874 15328
rect 17840 15287 17874 15310
rect 17840 15269 17848 15287
rect 17866 15269 17874 15287
rect 17840 15254 17874 15269
rect 17797 15209 17849 15217
rect 17797 15191 17812 15209
rect 17830 15191 17849 15209
rect 17797 15182 17849 15191
rect 17959 15155 17993 15161
rect 17959 15137 17967 15155
rect 17985 15137 17993 15155
rect 17959 15132 17993 15137
rect 17805 15016 17839 15025
rect 17805 14998 17813 15016
rect 17831 14998 17839 15016
rect 17805 14989 17839 14998
rect 17769 14956 17803 14972
rect 17565 14938 17573 14956
rect 17591 14938 17654 14956
rect 17565 14907 17599 14938
rect 17565 14889 17573 14907
rect 17591 14889 17600 14907
rect 17565 14874 17599 14889
rect 17501 14834 17519 14874
rect 17315 14817 17349 14826
rect 17315 14799 17323 14817
rect 17341 14799 17349 14817
rect 17315 14790 17349 14799
rect 17385 14816 17519 14834
rect 17385 14774 17403 14816
rect 17501 14775 17519 14816
rect 17555 14819 17590 14828
rect 17555 14801 17562 14819
rect 17580 14801 17590 14819
rect 17636 14819 17654 14938
rect 17732 14938 17777 14956
rect 17795 14938 17803 14956
rect 17732 14912 17750 14938
rect 17713 14906 17750 14912
rect 17769 14906 17803 14938
rect 17713 14888 17716 14906
rect 17734 14889 17750 14906
rect 17734 14888 17738 14889
rect 17767 14888 17777 14906
rect 17795 14888 17803 14906
rect 17713 14881 17738 14888
rect 17769 14873 17803 14888
rect 17841 14955 17875 14972
rect 17841 14937 17849 14955
rect 17867 14937 17875 14955
rect 17841 14906 17875 14937
rect 17841 14888 17849 14906
rect 17867 14888 17875 14906
rect 17841 14873 17875 14888
rect 17849 14830 17867 14873
rect 17965 14830 17983 15132
rect 17779 14819 17813 14828
rect 17636 14801 17787 14819
rect 17805 14801 17813 14819
rect 17555 14792 17590 14801
rect 17779 14792 17813 14801
rect 17849 14812 17983 14830
rect 17305 14765 17339 14773
rect 17305 14747 17313 14765
rect 17331 14747 17339 14765
rect 17305 14727 17339 14747
rect 17305 14709 17313 14727
rect 17331 14709 17339 14727
rect 17305 14689 17339 14709
rect 17305 14671 17313 14689
rect 17331 14671 17339 14689
rect 17305 14650 17339 14671
rect 17305 14632 17313 14650
rect 17331 14632 17339 14650
rect 17305 14609 17339 14632
rect 17305 14591 17313 14609
rect 17331 14591 17339 14609
rect 17305 14576 17339 14591
rect 17377 14765 17411 14774
rect 17377 14747 17385 14765
rect 17403 14747 17411 14765
rect 17377 14727 17411 14747
rect 17377 14709 17385 14727
rect 17403 14709 17411 14727
rect 17377 14689 17411 14709
rect 17377 14671 17385 14689
rect 17403 14671 17411 14689
rect 17493 14759 17527 14775
rect 17493 14741 17501 14759
rect 17519 14741 17527 14759
rect 17493 14709 17527 14741
rect 17493 14691 17501 14709
rect 17519 14691 17527 14709
rect 17493 14676 17527 14691
rect 17565 14758 17599 14775
rect 17849 14774 17867 14812
rect 17565 14740 17573 14758
rect 17591 14740 17599 14758
rect 17565 14709 17599 14740
rect 17565 14691 17573 14709
rect 17591 14691 17599 14709
rect 17565 14676 17599 14691
rect 17769 14758 17803 14774
rect 17769 14740 17777 14758
rect 17795 14740 17803 14758
rect 17769 14708 17803 14740
rect 17769 14690 17777 14708
rect 17795 14690 17803 14708
rect 17377 14650 17411 14671
rect 17377 14632 17385 14650
rect 17403 14632 17411 14650
rect 17377 14609 17411 14632
rect 17377 14591 17385 14609
rect 17403 14591 17411 14609
rect 17377 14576 17411 14591
rect 17313 14506 17331 14576
rect 17573 14506 17591 14676
rect 17769 14675 17803 14690
rect 17841 14757 17875 14774
rect 17965 14773 17983 14812
rect 18019 14818 18053 14827
rect 18019 14800 18027 14818
rect 18045 14800 18053 14818
rect 18019 14791 18053 14800
rect 17841 14739 17849 14757
rect 17867 14739 17875 14757
rect 17841 14708 17875 14739
rect 17841 14690 17849 14708
rect 17867 14690 17875 14708
rect 17841 14675 17875 14690
rect 17957 14765 17991 14773
rect 17957 14747 17965 14765
rect 17983 14747 17991 14765
rect 17957 14727 17991 14747
rect 17957 14709 17965 14727
rect 17983 14709 17991 14727
rect 17957 14689 17991 14709
rect 17777 14506 17795 14675
rect 17957 14671 17965 14689
rect 17983 14671 17991 14689
rect 17957 14650 17991 14671
rect 17957 14632 17965 14650
rect 17983 14632 17991 14650
rect 17957 14609 17991 14632
rect 17957 14591 17965 14609
rect 17983 14591 17991 14609
rect 17957 14576 17991 14591
rect 18029 14765 18063 14774
rect 18029 14747 18037 14765
rect 18055 14747 18063 14765
rect 18029 14727 18063 14747
rect 18029 14709 18037 14727
rect 18055 14709 18063 14727
rect 18029 14689 18063 14709
rect 18029 14671 18037 14689
rect 18055 14671 18063 14689
rect 18029 14650 18063 14671
rect 18029 14632 18037 14650
rect 18055 14632 18063 14650
rect 18029 14609 18063 14632
rect 18029 14591 18037 14609
rect 18055 14591 18063 14609
rect 18029 14576 18063 14591
rect 18037 14506 18055 14576
rect 17297 14500 18057 14506
rect 17297 14482 17313 14500
rect 17331 14482 17366 14500
rect 17384 14482 17417 14500
rect 17435 14482 17463 14500
rect 17481 14482 17509 14500
rect 17527 14482 17553 14500
rect 17571 14482 17601 14500
rect 17619 14482 17654 14500
rect 17672 14482 17705 14500
rect 17723 14482 17751 14500
rect 17769 14482 17797 14500
rect 17815 14482 17841 14500
rect 17859 14482 17884 14500
rect 17902 14482 17926 14500
rect 17944 14482 17966 14500
rect 17984 14482 18003 14500
rect 18021 14482 18034 14500
rect 18052 14482 18057 14500
rect 17297 14475 18057 14482
rect 18209 14344 18241 15566
rect 18670 15404 18702 15566
rect 18670 15402 18908 15404
rect 18670 15401 19305 15402
rect 18670 15398 19324 15401
rect 19431 15398 19462 15924
rect 19669 15843 19689 15924
rect 19935 15871 19954 15924
rect 20205 15871 20224 15925
rect 20355 15924 20496 15925
rect 19934 15845 19954 15871
rect 20204 15845 20224 15871
rect 18670 15396 19462 15398
rect 18670 15378 18880 15396
rect 18898 15378 18926 15396
rect 18944 15378 18980 15396
rect 18998 15378 19033 15396
rect 19051 15378 19084 15396
rect 19102 15378 19130 15396
rect 19148 15378 19176 15396
rect 19194 15378 19220 15396
rect 19238 15378 19263 15396
rect 19281 15378 19462 15396
rect 18670 15376 19462 15378
rect 19662 15828 19696 15843
rect 19662 15810 19670 15828
rect 19688 15810 19696 15828
rect 19662 15787 19696 15810
rect 19662 15769 19670 15787
rect 19688 15769 19696 15787
rect 19662 15748 19696 15769
rect 19662 15730 19670 15748
rect 19688 15730 19696 15748
rect 19662 15710 19696 15730
rect 19662 15692 19670 15710
rect 19688 15692 19696 15710
rect 19662 15672 19696 15692
rect 19662 15654 19670 15672
rect 19688 15654 19696 15672
rect 19662 15628 19696 15654
rect 19662 15610 19670 15628
rect 19688 15610 19696 15628
rect 19662 15587 19696 15610
rect 19662 15569 19670 15587
rect 19688 15569 19696 15587
rect 19662 15548 19696 15569
rect 19662 15530 19670 15548
rect 19688 15530 19696 15548
rect 19662 15510 19696 15530
rect 19662 15492 19670 15510
rect 19688 15492 19696 15510
rect 19662 15472 19696 15492
rect 19662 15454 19670 15472
rect 19688 15454 19696 15472
rect 19662 15428 19696 15454
rect 19662 15410 19670 15428
rect 19688 15410 19696 15428
rect 19662 15387 19696 15410
rect 18670 15372 19461 15376
rect 18838 15371 19324 15372
rect 18838 15370 18870 15371
rect 18838 15309 18856 15370
rect 18839 15307 18856 15309
rect 18839 15288 18857 15307
rect 18831 15273 18865 15288
rect 18831 15255 18839 15273
rect 18857 15255 18865 15273
rect 18831 15232 18865 15255
rect 18831 15214 18839 15232
rect 18857 15214 18865 15232
rect 18831 15193 18865 15214
rect 18831 15175 18839 15193
rect 18857 15175 18865 15193
rect 18831 15155 18865 15175
rect 18831 15137 18839 15155
rect 18857 15137 18865 15155
rect 18831 15117 18865 15137
rect 18831 15099 18839 15117
rect 18857 15099 18865 15117
rect 18831 15091 18865 15099
rect 18903 15273 18937 15288
rect 19269 15286 19287 15371
rect 19662 15369 19670 15387
rect 19688 15369 19696 15387
rect 19662 15348 19696 15369
rect 19662 15330 19670 15348
rect 19688 15330 19696 15348
rect 19662 15310 19696 15330
rect 19662 15292 19670 15310
rect 19688 15292 19696 15310
rect 18903 15255 18911 15273
rect 18929 15255 18937 15273
rect 18903 15232 18937 15255
rect 18903 15214 18911 15232
rect 18929 15214 18937 15232
rect 18903 15193 18937 15214
rect 18903 15175 18911 15193
rect 18929 15175 18937 15193
rect 18903 15155 18937 15175
rect 18903 15137 18911 15155
rect 18929 15137 18937 15155
rect 18903 15117 18937 15137
rect 18903 15099 18911 15117
rect 18929 15099 18937 15117
rect 18903 15090 18937 15099
rect 19261 15271 19295 15286
rect 19261 15253 19269 15271
rect 19287 15253 19295 15271
rect 19261 15230 19295 15253
rect 19261 15212 19269 15230
rect 19287 15212 19295 15230
rect 19261 15191 19295 15212
rect 19261 15173 19269 15191
rect 19287 15173 19295 15191
rect 19261 15153 19295 15173
rect 19261 15135 19269 15153
rect 19287 15135 19295 15153
rect 19261 15115 19295 15135
rect 19261 15097 19269 15115
rect 19287 15097 19295 15115
rect 18911 15086 18929 15090
rect 19261 15089 19295 15097
rect 19333 15271 19367 15286
rect 19333 15253 19341 15271
rect 19359 15253 19367 15271
rect 19333 15230 19367 15253
rect 19333 15212 19341 15230
rect 19359 15212 19367 15230
rect 19333 15191 19367 15212
rect 19333 15173 19341 15191
rect 19359 15173 19367 15191
rect 19333 15153 19367 15173
rect 19333 15135 19341 15153
rect 19359 15135 19367 15153
rect 19333 15115 19367 15135
rect 19333 15097 19341 15115
rect 19359 15097 19367 15115
rect 19333 15088 19367 15097
rect 19662 15272 19696 15292
rect 19662 15254 19670 15272
rect 19688 15254 19696 15272
rect 19662 15228 19696 15254
rect 19662 15210 19670 15228
rect 19688 15210 19696 15228
rect 19662 15187 19696 15210
rect 19662 15169 19670 15187
rect 19688 15169 19696 15187
rect 19662 15148 19696 15169
rect 19662 15130 19670 15148
rect 19688 15130 19696 15148
rect 19662 15110 19696 15130
rect 19662 15092 19670 15110
rect 19688 15092 19696 15110
rect 18841 15069 18875 15074
rect 18726 15065 18875 15069
rect 18726 15047 18849 15065
rect 18867 15047 18875 15065
rect 18726 15045 18875 15047
rect 18271 15019 18305 15028
rect 18271 15001 18279 15019
rect 18297 15001 18305 15019
rect 18271 14992 18305 15001
rect 18330 14824 18361 14836
rect 18322 14817 18361 14824
rect 18322 14800 18337 14817
rect 18354 14800 18361 14817
rect 18322 14790 18361 14800
rect 18330 14780 18361 14790
rect 17161 14338 18241 14344
rect 17161 14320 17277 14338
rect 17295 14320 17323 14338
rect 17341 14320 17377 14338
rect 17395 14320 17430 14338
rect 17448 14320 17481 14338
rect 17499 14320 17527 14338
rect 17545 14320 17573 14338
rect 17591 14320 17617 14338
rect 17635 14320 17660 14338
rect 17678 14320 17704 14338
rect 17722 14320 17750 14338
rect 17768 14320 17804 14338
rect 17822 14320 17857 14338
rect 17875 14320 17908 14338
rect 17926 14320 17954 14338
rect 17972 14320 18000 14338
rect 18018 14320 18044 14338
rect 18062 14320 18087 14338
rect 18105 14320 18241 14338
rect 17161 14313 18241 14320
rect 17361 14234 17379 14313
rect 17353 14226 17387 14234
rect 17353 14208 17361 14226
rect 17379 14208 17387 14226
rect 17353 14188 17387 14208
rect 17353 14170 17361 14188
rect 17379 14170 17387 14188
rect 17353 14150 17387 14170
rect 17353 14132 17361 14150
rect 17379 14132 17387 14150
rect 17353 14111 17387 14132
rect 17353 14093 17361 14111
rect 17379 14093 17387 14111
rect 17353 14070 17387 14093
rect 17353 14052 17361 14070
rect 17379 14052 17387 14070
rect 17353 14037 17387 14052
rect 17425 14226 17459 14235
rect 17982 14233 18000 14313
rect 18112 14312 18241 14313
rect 18342 14760 18361 14780
rect 17425 14208 17433 14226
rect 17451 14208 17459 14226
rect 17425 14188 17459 14208
rect 17425 14170 17433 14188
rect 17451 14170 17459 14188
rect 17425 14150 17459 14170
rect 17425 14132 17433 14150
rect 17451 14132 17459 14150
rect 17425 14111 17459 14132
rect 17425 14093 17433 14111
rect 17451 14093 17459 14111
rect 17425 14070 17459 14093
rect 17425 14052 17433 14070
rect 17451 14052 17459 14070
rect 17425 14037 17459 14052
rect 17903 14224 17936 14232
rect 17903 14206 17910 14224
rect 17928 14206 17936 14224
rect 17903 14186 17936 14206
rect 17903 14168 17910 14186
rect 17928 14168 17936 14186
rect 17903 14148 17936 14168
rect 17903 14130 17910 14148
rect 17928 14130 17936 14148
rect 17903 14109 17936 14130
rect 17903 14091 17910 14109
rect 17928 14091 17936 14109
rect 17903 14068 17936 14091
rect 17903 14050 17910 14068
rect 17928 14050 17936 14068
rect 17363 13998 17397 14007
rect 17363 13980 17371 13998
rect 17389 13980 17397 13998
rect 17363 13971 17397 13980
rect 17430 13949 17453 14037
rect 17903 14035 17936 14050
rect 17974 14224 18008 14233
rect 17974 14206 17982 14224
rect 18000 14206 18008 14224
rect 17974 14186 18008 14206
rect 17974 14168 17982 14186
rect 18000 14168 18008 14186
rect 17974 14148 18008 14168
rect 17974 14130 17982 14148
rect 18000 14130 18008 14148
rect 17974 14109 18008 14130
rect 17974 14091 17982 14109
rect 18000 14091 18008 14109
rect 17974 14068 18008 14091
rect 17974 14050 17982 14068
rect 18000 14050 18008 14068
rect 17974 14035 18008 14050
rect 17045 13931 17453 13949
rect 17363 13876 17397 13885
rect 16256 13858 17371 13876
rect 17389 13858 17397 13876
rect 17363 13849 17397 13858
rect 17430 13832 17453 13931
rect 17908 13949 17929 14035
rect 17964 13994 17998 14003
rect 17964 13976 17972 13994
rect 17990 13976 17998 13994
rect 17964 13967 17998 13976
rect 18342 13949 18360 14760
rect 18726 14430 18750 15045
rect 18841 15038 18875 15045
rect 18912 15064 18929 15086
rect 19341 15084 19359 15088
rect 19271 15067 19305 15072
rect 19156 15064 19305 15067
rect 18912 15063 19305 15064
rect 18912 15045 19279 15063
rect 19297 15045 19305 15063
rect 18912 15043 19305 15045
rect 18912 15040 19180 15043
rect 18912 15030 18930 15040
rect 18913 15023 18930 15030
rect 18843 14975 18877 14984
rect 18843 14957 18851 14975
rect 18869 14957 18877 14975
rect 18843 14948 18877 14957
rect 18913 14932 18931 15023
rect 18833 14923 18867 14931
rect 18833 14905 18841 14923
rect 18859 14905 18867 14923
rect 18833 14885 18867 14905
rect 18833 14867 18841 14885
rect 18859 14867 18867 14885
rect 18833 14847 18867 14867
rect 18833 14829 18841 14847
rect 18859 14829 18867 14847
rect 18833 14808 18867 14829
rect 18833 14790 18841 14808
rect 18859 14790 18867 14808
rect 18833 14767 18867 14790
rect 18833 14749 18841 14767
rect 18859 14749 18867 14767
rect 18833 14734 18867 14749
rect 18905 14923 18939 14932
rect 18905 14905 18913 14923
rect 18931 14905 18939 14923
rect 18905 14885 18939 14905
rect 18905 14867 18913 14885
rect 18931 14867 18939 14885
rect 18905 14847 18939 14867
rect 18905 14829 18913 14847
rect 18931 14829 18939 14847
rect 18905 14808 18939 14829
rect 18905 14790 18913 14808
rect 18931 14790 18939 14808
rect 18905 14767 18939 14790
rect 18905 14749 18913 14767
rect 18931 14749 18939 14767
rect 18905 14734 18939 14749
rect 18841 14650 18859 14734
rect 18833 14635 18867 14650
rect 18833 14617 18841 14635
rect 18859 14617 18867 14635
rect 18833 14594 18867 14617
rect 18833 14576 18841 14594
rect 18859 14576 18867 14594
rect 18833 14555 18867 14576
rect 18833 14537 18841 14555
rect 18859 14537 18867 14555
rect 18833 14517 18867 14537
rect 18833 14499 18841 14517
rect 18859 14499 18867 14517
rect 18833 14479 18867 14499
rect 18833 14461 18841 14479
rect 18859 14461 18867 14479
rect 18833 14453 18867 14461
rect 18905 14635 18939 14650
rect 18905 14617 18913 14635
rect 18931 14617 18939 14635
rect 18905 14594 18939 14617
rect 18905 14576 18913 14594
rect 18931 14576 18939 14594
rect 18905 14555 18939 14576
rect 18905 14537 18913 14555
rect 18931 14537 18939 14555
rect 18905 14517 18939 14537
rect 18905 14499 18913 14517
rect 18931 14499 18939 14517
rect 18905 14479 18939 14499
rect 18905 14461 18913 14479
rect 18931 14461 18939 14479
rect 18905 14452 18939 14461
rect 18843 14430 18877 14436
rect 18726 14427 18877 14430
rect 18726 14409 18851 14427
rect 18869 14409 18877 14427
rect 18726 14406 18877 14409
rect 18843 14400 18877 14406
rect 18913 14410 18931 14452
rect 19156 14428 19180 15040
rect 19271 15036 19305 15043
rect 19342 15046 19359 15084
rect 19662 15072 19696 15092
rect 19662 15054 19670 15072
rect 19688 15054 19696 15072
rect 19662 15046 19696 15054
rect 19734 15828 19768 15843
rect 19734 15810 19742 15828
rect 19760 15810 19768 15828
rect 19734 15787 19768 15810
rect 19734 15769 19742 15787
rect 19760 15769 19768 15787
rect 19734 15748 19768 15769
rect 19734 15730 19742 15748
rect 19760 15730 19768 15748
rect 19734 15710 19768 15730
rect 19734 15692 19742 15710
rect 19760 15692 19768 15710
rect 19734 15672 19768 15692
rect 19734 15654 19742 15672
rect 19760 15654 19768 15672
rect 19734 15628 19768 15654
rect 19734 15610 19742 15628
rect 19760 15610 19768 15628
rect 19734 15587 19768 15610
rect 19734 15569 19742 15587
rect 19760 15569 19768 15587
rect 19734 15548 19768 15569
rect 19734 15530 19742 15548
rect 19760 15530 19768 15548
rect 19734 15510 19768 15530
rect 19734 15492 19742 15510
rect 19760 15492 19768 15510
rect 19734 15472 19768 15492
rect 19734 15454 19742 15472
rect 19760 15454 19768 15472
rect 19734 15428 19768 15454
rect 19734 15410 19742 15428
rect 19760 15410 19768 15428
rect 19734 15387 19768 15410
rect 19734 15369 19742 15387
rect 19760 15369 19768 15387
rect 19734 15348 19768 15369
rect 19734 15330 19742 15348
rect 19760 15330 19768 15348
rect 19734 15310 19768 15330
rect 19734 15292 19742 15310
rect 19760 15292 19768 15310
rect 19734 15272 19768 15292
rect 19734 15254 19742 15272
rect 19760 15254 19768 15272
rect 19734 15228 19768 15254
rect 19734 15210 19742 15228
rect 19760 15210 19768 15228
rect 19734 15187 19768 15210
rect 19734 15169 19742 15187
rect 19760 15169 19768 15187
rect 19734 15148 19768 15169
rect 19734 15130 19742 15148
rect 19760 15130 19768 15148
rect 19734 15110 19768 15130
rect 19734 15092 19742 15110
rect 19760 15092 19768 15110
rect 19734 15072 19768 15092
rect 19734 15054 19742 15072
rect 19760 15054 19768 15072
rect 19342 15028 19360 15046
rect 19734 15045 19768 15054
rect 19927 15830 19961 15845
rect 19927 15812 19935 15830
rect 19953 15812 19961 15830
rect 19927 15789 19961 15812
rect 19927 15771 19935 15789
rect 19953 15771 19961 15789
rect 19927 15750 19961 15771
rect 19927 15732 19935 15750
rect 19953 15732 19961 15750
rect 19927 15712 19961 15732
rect 19927 15694 19935 15712
rect 19953 15694 19961 15712
rect 19927 15674 19961 15694
rect 19927 15656 19935 15674
rect 19953 15656 19961 15674
rect 19927 15630 19961 15656
rect 19927 15612 19935 15630
rect 19953 15612 19961 15630
rect 19927 15589 19961 15612
rect 19927 15571 19935 15589
rect 19953 15571 19961 15589
rect 19927 15550 19961 15571
rect 19927 15532 19935 15550
rect 19953 15532 19961 15550
rect 19927 15512 19961 15532
rect 19927 15494 19935 15512
rect 19953 15494 19961 15512
rect 19927 15474 19961 15494
rect 19927 15456 19935 15474
rect 19953 15456 19961 15474
rect 19927 15430 19961 15456
rect 19927 15412 19935 15430
rect 19953 15412 19961 15430
rect 19927 15389 19961 15412
rect 19927 15371 19935 15389
rect 19953 15371 19961 15389
rect 19927 15350 19961 15371
rect 19927 15332 19935 15350
rect 19953 15332 19961 15350
rect 19927 15312 19961 15332
rect 19927 15294 19935 15312
rect 19953 15294 19961 15312
rect 19927 15274 19961 15294
rect 19927 15256 19935 15274
rect 19953 15256 19961 15274
rect 19927 15230 19961 15256
rect 19927 15212 19935 15230
rect 19953 15212 19961 15230
rect 19927 15189 19961 15212
rect 19927 15171 19935 15189
rect 19953 15171 19961 15189
rect 19927 15150 19961 15171
rect 19927 15132 19935 15150
rect 19953 15132 19961 15150
rect 19927 15112 19961 15132
rect 19927 15094 19935 15112
rect 19953 15094 19961 15112
rect 19927 15074 19961 15094
rect 19927 15056 19935 15074
rect 19953 15056 19961 15074
rect 19927 15048 19961 15056
rect 19999 15830 20033 15845
rect 19999 15812 20007 15830
rect 20025 15812 20033 15830
rect 19999 15789 20033 15812
rect 19999 15771 20007 15789
rect 20025 15771 20033 15789
rect 19999 15750 20033 15771
rect 19999 15732 20007 15750
rect 20025 15732 20033 15750
rect 19999 15712 20033 15732
rect 19999 15694 20007 15712
rect 20025 15694 20033 15712
rect 19999 15674 20033 15694
rect 19999 15656 20007 15674
rect 20025 15656 20033 15674
rect 19999 15630 20033 15656
rect 19999 15612 20007 15630
rect 20025 15612 20033 15630
rect 19999 15589 20033 15612
rect 19999 15571 20007 15589
rect 20025 15571 20033 15589
rect 19999 15550 20033 15571
rect 19999 15532 20007 15550
rect 20025 15532 20033 15550
rect 19999 15512 20033 15532
rect 19999 15494 20007 15512
rect 20025 15494 20033 15512
rect 19999 15474 20033 15494
rect 19999 15456 20007 15474
rect 20025 15456 20033 15474
rect 19999 15430 20033 15456
rect 19999 15412 20007 15430
rect 20025 15412 20033 15430
rect 19999 15389 20033 15412
rect 19999 15371 20007 15389
rect 20025 15371 20033 15389
rect 19999 15350 20033 15371
rect 19999 15332 20007 15350
rect 20025 15332 20033 15350
rect 19999 15312 20033 15332
rect 19999 15294 20007 15312
rect 20025 15294 20033 15312
rect 19999 15274 20033 15294
rect 19999 15256 20007 15274
rect 20025 15256 20033 15274
rect 19999 15230 20033 15256
rect 19999 15212 20007 15230
rect 20025 15212 20033 15230
rect 19999 15189 20033 15212
rect 19999 15171 20007 15189
rect 20025 15171 20033 15189
rect 19999 15150 20033 15171
rect 19999 15132 20007 15150
rect 20025 15132 20033 15150
rect 19999 15112 20033 15132
rect 19999 15094 20007 15112
rect 20025 15094 20033 15112
rect 19999 15074 20033 15094
rect 19999 15056 20007 15074
rect 20025 15056 20033 15074
rect 19999 15047 20033 15056
rect 20197 15830 20231 15845
rect 20197 15812 20205 15830
rect 20223 15812 20231 15830
rect 20197 15789 20231 15812
rect 20197 15771 20205 15789
rect 20223 15771 20231 15789
rect 20197 15750 20231 15771
rect 20197 15732 20205 15750
rect 20223 15732 20231 15750
rect 20197 15712 20231 15732
rect 20197 15694 20205 15712
rect 20223 15694 20231 15712
rect 20197 15674 20231 15694
rect 20197 15656 20205 15674
rect 20223 15656 20231 15674
rect 20197 15630 20231 15656
rect 20197 15612 20205 15630
rect 20223 15612 20231 15630
rect 20197 15589 20231 15612
rect 20197 15571 20205 15589
rect 20223 15571 20231 15589
rect 20197 15550 20231 15571
rect 20197 15532 20205 15550
rect 20223 15532 20231 15550
rect 20197 15512 20231 15532
rect 20197 15494 20205 15512
rect 20223 15494 20231 15512
rect 20197 15474 20231 15494
rect 20197 15456 20205 15474
rect 20223 15456 20231 15474
rect 20197 15430 20231 15456
rect 20197 15412 20205 15430
rect 20223 15412 20231 15430
rect 20197 15389 20231 15412
rect 20197 15371 20205 15389
rect 20223 15371 20231 15389
rect 20197 15350 20231 15371
rect 20197 15332 20205 15350
rect 20223 15332 20231 15350
rect 20197 15312 20231 15332
rect 20197 15294 20205 15312
rect 20223 15294 20231 15312
rect 20197 15274 20231 15294
rect 20197 15256 20205 15274
rect 20223 15256 20231 15274
rect 20197 15230 20231 15256
rect 20197 15212 20205 15230
rect 20223 15212 20231 15230
rect 20197 15189 20231 15212
rect 20197 15171 20205 15189
rect 20223 15171 20231 15189
rect 20197 15150 20231 15171
rect 20197 15132 20205 15150
rect 20223 15132 20231 15150
rect 20197 15112 20231 15132
rect 20197 15094 20205 15112
rect 20223 15094 20231 15112
rect 20197 15074 20231 15094
rect 20197 15056 20205 15074
rect 20223 15056 20231 15074
rect 20197 15048 20231 15056
rect 20269 15830 20303 15845
rect 20475 15843 20495 15924
rect 20269 15812 20277 15830
rect 20295 15812 20303 15830
rect 20269 15789 20303 15812
rect 20269 15771 20277 15789
rect 20295 15771 20303 15789
rect 20269 15750 20303 15771
rect 20269 15732 20277 15750
rect 20295 15732 20303 15750
rect 20269 15712 20303 15732
rect 20269 15694 20277 15712
rect 20295 15694 20303 15712
rect 20269 15674 20303 15694
rect 20269 15656 20277 15674
rect 20295 15656 20303 15674
rect 20269 15630 20303 15656
rect 20269 15612 20277 15630
rect 20295 15612 20303 15630
rect 20269 15589 20303 15612
rect 20269 15571 20277 15589
rect 20295 15571 20303 15589
rect 20269 15550 20303 15571
rect 20269 15532 20277 15550
rect 20295 15532 20303 15550
rect 20269 15512 20303 15532
rect 20269 15494 20277 15512
rect 20295 15494 20303 15512
rect 20269 15474 20303 15494
rect 20269 15456 20277 15474
rect 20295 15456 20303 15474
rect 20269 15430 20303 15456
rect 20269 15412 20277 15430
rect 20295 15412 20303 15430
rect 20269 15389 20303 15412
rect 20269 15371 20277 15389
rect 20295 15371 20303 15389
rect 20269 15350 20303 15371
rect 20269 15332 20277 15350
rect 20295 15332 20303 15350
rect 20269 15312 20303 15332
rect 20269 15294 20277 15312
rect 20295 15294 20303 15312
rect 20269 15274 20303 15294
rect 20269 15256 20277 15274
rect 20295 15256 20303 15274
rect 20269 15230 20303 15256
rect 20269 15212 20277 15230
rect 20295 15212 20303 15230
rect 20269 15189 20303 15212
rect 20269 15171 20277 15189
rect 20295 15171 20303 15189
rect 20269 15150 20303 15171
rect 20269 15132 20277 15150
rect 20295 15132 20303 15150
rect 20269 15112 20303 15132
rect 20269 15094 20277 15112
rect 20295 15094 20303 15112
rect 20269 15074 20303 15094
rect 20269 15056 20277 15074
rect 20295 15056 20303 15074
rect 20269 15047 20303 15056
rect 20468 15828 20502 15843
rect 20468 15810 20476 15828
rect 20494 15810 20502 15828
rect 20468 15787 20502 15810
rect 20468 15769 20476 15787
rect 20494 15769 20502 15787
rect 20468 15748 20502 15769
rect 20468 15730 20476 15748
rect 20494 15730 20502 15748
rect 20468 15710 20502 15730
rect 20468 15692 20476 15710
rect 20494 15692 20502 15710
rect 20468 15672 20502 15692
rect 20468 15654 20476 15672
rect 20494 15654 20502 15672
rect 20468 15628 20502 15654
rect 20468 15610 20476 15628
rect 20494 15610 20502 15628
rect 20468 15587 20502 15610
rect 20468 15569 20476 15587
rect 20494 15569 20502 15587
rect 20468 15548 20502 15569
rect 20468 15530 20476 15548
rect 20494 15530 20502 15548
rect 20468 15510 20502 15530
rect 20468 15492 20476 15510
rect 20494 15492 20502 15510
rect 20468 15472 20502 15492
rect 20468 15454 20476 15472
rect 20494 15454 20502 15472
rect 20468 15428 20502 15454
rect 20468 15410 20476 15428
rect 20494 15410 20502 15428
rect 20468 15387 20502 15410
rect 20468 15369 20476 15387
rect 20494 15369 20502 15387
rect 20468 15348 20502 15369
rect 20468 15330 20476 15348
rect 20494 15330 20502 15348
rect 20468 15310 20502 15330
rect 20468 15292 20476 15310
rect 20494 15292 20502 15310
rect 20468 15272 20502 15292
rect 20468 15254 20476 15272
rect 20494 15254 20502 15272
rect 20468 15228 20502 15254
rect 20468 15210 20476 15228
rect 20494 15210 20502 15228
rect 20468 15187 20502 15210
rect 20468 15169 20476 15187
rect 20494 15169 20502 15187
rect 20468 15148 20502 15169
rect 20468 15130 20476 15148
rect 20494 15130 20502 15148
rect 20468 15110 20502 15130
rect 20468 15092 20476 15110
rect 20494 15092 20502 15110
rect 20468 15072 20502 15092
rect 20468 15054 20476 15072
rect 20494 15054 20502 15072
rect 19742 15041 19760 15045
rect 20007 15043 20025 15047
rect 20277 15043 20295 15047
rect 20468 15046 20502 15054
rect 20540 15828 20574 15843
rect 20540 15810 20548 15828
rect 20566 15810 20574 15828
rect 20540 15787 20574 15810
rect 20540 15769 20548 15787
rect 20566 15769 20574 15787
rect 20540 15748 20574 15769
rect 20540 15730 20548 15748
rect 20566 15730 20574 15748
rect 20540 15710 20574 15730
rect 20540 15692 20548 15710
rect 20566 15692 20574 15710
rect 20540 15672 20574 15692
rect 20540 15654 20548 15672
rect 20566 15654 20574 15672
rect 20540 15628 20574 15654
rect 20540 15610 20548 15628
rect 20566 15610 20574 15628
rect 20540 15587 20574 15610
rect 20540 15569 20548 15587
rect 20566 15569 20574 15587
rect 20540 15548 20574 15569
rect 20540 15530 20548 15548
rect 20566 15530 20574 15548
rect 20540 15510 20574 15530
rect 20540 15492 20548 15510
rect 20566 15492 20574 15510
rect 20540 15472 20574 15492
rect 20540 15454 20548 15472
rect 20566 15454 20574 15472
rect 20540 15428 20574 15454
rect 20540 15410 20548 15428
rect 20566 15410 20574 15428
rect 20540 15387 20574 15410
rect 20540 15369 20548 15387
rect 20566 15369 20574 15387
rect 20540 15348 20574 15369
rect 20540 15330 20548 15348
rect 20566 15330 20574 15348
rect 20540 15310 20574 15330
rect 20540 15292 20548 15310
rect 20566 15292 20574 15310
rect 20540 15272 20574 15292
rect 20540 15254 20548 15272
rect 20566 15254 20574 15272
rect 20540 15228 20574 15254
rect 20540 15210 20548 15228
rect 20566 15210 20574 15228
rect 20540 15187 20574 15210
rect 20540 15169 20548 15187
rect 20566 15169 20574 15187
rect 20540 15148 20574 15169
rect 20540 15130 20548 15148
rect 20566 15130 20574 15148
rect 20540 15110 20574 15130
rect 20540 15092 20548 15110
rect 20566 15092 20574 15110
rect 20540 15072 20574 15092
rect 20540 15054 20548 15072
rect 20566 15054 20574 15072
rect 20540 15045 20574 15054
rect 19343 15021 19360 15028
rect 19343 14990 19361 15021
rect 19743 15016 19760 15041
rect 20008 15018 20025 15043
rect 20278 15018 20295 15043
rect 20548 15041 20566 15045
rect 19672 14993 19706 14998
rect 19635 14990 19706 14993
rect 19343 14989 19706 14990
rect 19273 14973 19307 14982
rect 19273 14955 19281 14973
rect 19299 14955 19307 14973
rect 19273 14946 19307 14955
rect 19343 14972 19680 14989
rect 19343 14930 19361 14972
rect 19635 14971 19680 14972
rect 19698 14971 19706 14989
rect 19635 14969 19706 14971
rect 19672 14962 19706 14969
rect 19742 14993 19760 15016
rect 19937 14995 19971 15000
rect 19900 14993 19971 14995
rect 19742 14991 19971 14993
rect 19742 14975 19945 14991
rect 19263 14921 19297 14929
rect 19263 14903 19271 14921
rect 19289 14903 19297 14921
rect 19263 14883 19297 14903
rect 19263 14865 19271 14883
rect 19289 14865 19297 14883
rect 19263 14845 19297 14865
rect 19263 14827 19271 14845
rect 19289 14827 19297 14845
rect 19263 14806 19297 14827
rect 19263 14788 19271 14806
rect 19289 14788 19297 14806
rect 19263 14765 19297 14788
rect 19263 14747 19271 14765
rect 19289 14747 19297 14765
rect 19263 14732 19297 14747
rect 19335 14921 19369 14930
rect 19742 14929 19760 14975
rect 19899 14973 19945 14975
rect 19963 14973 19971 14991
rect 19899 14971 19971 14973
rect 19937 14964 19971 14971
rect 20007 14989 20025 15018
rect 20207 14995 20241 15000
rect 20170 14991 20241 14995
rect 20170 14989 20215 14991
rect 20007 14973 20215 14989
rect 20233 14973 20241 14991
rect 20007 14971 20241 14973
rect 20007 14931 20025 14971
rect 20170 14969 20241 14971
rect 20207 14964 20241 14969
rect 20277 14989 20295 15018
rect 20549 15016 20566 15041
rect 20478 14993 20512 14998
rect 20441 14989 20512 14993
rect 20277 14971 20486 14989
rect 20504 14971 20512 14989
rect 20277 14931 20295 14971
rect 20441 14969 20512 14971
rect 20478 14962 20512 14969
rect 20548 14987 20566 15016
rect 20631 14988 20665 14994
rect 20631 14987 20639 14988
rect 20548 14970 20639 14987
rect 20657 14987 20665 14988
rect 21811 14987 21829 16133
rect 22295 16095 22357 16133
rect 20657 14970 21829 14987
rect 20548 14969 21829 14970
rect 19335 14903 19343 14921
rect 19361 14903 19369 14921
rect 19335 14883 19369 14903
rect 19335 14865 19343 14883
rect 19361 14865 19369 14883
rect 19335 14845 19369 14865
rect 19335 14827 19343 14845
rect 19361 14827 19369 14845
rect 19335 14806 19369 14827
rect 19335 14788 19343 14806
rect 19361 14788 19369 14806
rect 19335 14765 19369 14788
rect 19335 14747 19343 14765
rect 19361 14747 19369 14765
rect 19335 14732 19369 14747
rect 19662 14920 19696 14928
rect 19662 14902 19670 14920
rect 19688 14902 19696 14920
rect 19662 14882 19696 14902
rect 19662 14864 19670 14882
rect 19688 14864 19696 14882
rect 19662 14844 19696 14864
rect 19662 14826 19670 14844
rect 19688 14826 19696 14844
rect 19662 14805 19696 14826
rect 19662 14787 19670 14805
rect 19688 14787 19696 14805
rect 19662 14764 19696 14787
rect 19662 14746 19670 14764
rect 19688 14746 19696 14764
rect 19271 14648 19289 14732
rect 19662 14731 19696 14746
rect 19734 14920 19768 14929
rect 19734 14902 19742 14920
rect 19760 14902 19768 14920
rect 19734 14882 19768 14902
rect 19734 14864 19742 14882
rect 19760 14864 19768 14882
rect 19734 14844 19768 14864
rect 19734 14826 19742 14844
rect 19760 14826 19768 14844
rect 19734 14805 19768 14826
rect 19734 14787 19742 14805
rect 19760 14787 19768 14805
rect 19734 14764 19768 14787
rect 19734 14746 19742 14764
rect 19760 14746 19768 14764
rect 19734 14731 19768 14746
rect 19927 14922 19961 14930
rect 19927 14904 19935 14922
rect 19953 14904 19961 14922
rect 19927 14884 19961 14904
rect 19927 14866 19935 14884
rect 19953 14866 19961 14884
rect 19927 14846 19961 14866
rect 19927 14828 19935 14846
rect 19953 14828 19961 14846
rect 19927 14807 19961 14828
rect 19927 14789 19935 14807
rect 19953 14789 19961 14807
rect 19927 14766 19961 14789
rect 19927 14748 19935 14766
rect 19953 14748 19961 14766
rect 19927 14733 19961 14748
rect 19999 14922 20033 14931
rect 19999 14904 20007 14922
rect 20025 14904 20033 14922
rect 19999 14884 20033 14904
rect 19999 14866 20007 14884
rect 20025 14866 20033 14884
rect 19999 14846 20033 14866
rect 19999 14828 20007 14846
rect 20025 14828 20033 14846
rect 19999 14807 20033 14828
rect 19999 14789 20007 14807
rect 20025 14789 20033 14807
rect 19999 14766 20033 14789
rect 19999 14748 20007 14766
rect 20025 14748 20033 14766
rect 19999 14733 20033 14748
rect 20197 14922 20231 14930
rect 20197 14904 20205 14922
rect 20223 14904 20231 14922
rect 20197 14884 20231 14904
rect 20197 14866 20205 14884
rect 20223 14866 20231 14884
rect 20197 14846 20231 14866
rect 20197 14828 20205 14846
rect 20223 14828 20231 14846
rect 20197 14807 20231 14828
rect 20197 14789 20205 14807
rect 20223 14789 20231 14807
rect 20197 14766 20231 14789
rect 20197 14748 20205 14766
rect 20223 14748 20231 14766
rect 20197 14733 20231 14748
rect 20269 14922 20303 14931
rect 20548 14929 20566 14969
rect 20631 14965 20665 14969
rect 20269 14904 20277 14922
rect 20295 14904 20303 14922
rect 20269 14884 20303 14904
rect 20269 14866 20277 14884
rect 20295 14866 20303 14884
rect 20269 14846 20303 14866
rect 20269 14828 20277 14846
rect 20295 14828 20303 14846
rect 20269 14807 20303 14828
rect 20269 14789 20277 14807
rect 20295 14789 20303 14807
rect 20269 14766 20303 14789
rect 20269 14748 20277 14766
rect 20295 14748 20303 14766
rect 20269 14733 20303 14748
rect 20468 14920 20502 14928
rect 20468 14902 20476 14920
rect 20494 14902 20502 14920
rect 20468 14882 20502 14902
rect 20468 14864 20476 14882
rect 20494 14864 20502 14882
rect 20468 14844 20502 14864
rect 20468 14826 20476 14844
rect 20494 14826 20502 14844
rect 20468 14805 20502 14826
rect 20468 14787 20476 14805
rect 20494 14787 20502 14805
rect 20468 14764 20502 14787
rect 20468 14746 20476 14764
rect 20494 14746 20502 14764
rect 19263 14633 19297 14648
rect 19263 14615 19271 14633
rect 19289 14615 19297 14633
rect 19263 14592 19297 14615
rect 19263 14574 19271 14592
rect 19289 14574 19297 14592
rect 19263 14553 19297 14574
rect 19263 14535 19271 14553
rect 19289 14535 19297 14553
rect 19263 14515 19297 14535
rect 19263 14497 19271 14515
rect 19289 14497 19297 14515
rect 19263 14477 19297 14497
rect 19263 14459 19271 14477
rect 19289 14459 19297 14477
rect 19263 14451 19297 14459
rect 19335 14633 19369 14648
rect 19335 14615 19343 14633
rect 19361 14615 19369 14633
rect 19670 14639 19688 14731
rect 19935 14643 19953 14733
rect 20205 14643 20223 14733
rect 20468 14731 20502 14746
rect 20540 14920 20574 14929
rect 20540 14902 20548 14920
rect 20566 14902 20574 14920
rect 20540 14882 20574 14902
rect 20540 14864 20548 14882
rect 20566 14864 20574 14882
rect 20540 14844 20574 14864
rect 20540 14826 20548 14844
rect 20566 14826 20574 14844
rect 20540 14805 20574 14826
rect 20540 14787 20548 14805
rect 20566 14787 20574 14805
rect 20540 14764 20574 14787
rect 20540 14746 20548 14764
rect 20566 14746 20574 14764
rect 20540 14731 20574 14746
rect 20476 14643 20494 14731
rect 19729 14639 20494 14643
rect 19670 14637 20494 14639
rect 19670 14621 19745 14637
rect 19335 14592 19369 14615
rect 19729 14619 19745 14621
rect 19763 14619 19798 14637
rect 19816 14619 19849 14637
rect 19867 14619 19895 14637
rect 19913 14619 19941 14637
rect 19959 14619 19985 14637
rect 20003 14619 20033 14637
rect 20051 14619 20086 14637
rect 20104 14619 20137 14637
rect 20155 14619 20183 14637
rect 20201 14619 20229 14637
rect 20247 14619 20273 14637
rect 20291 14619 20316 14637
rect 20334 14619 20358 14637
rect 20376 14619 20398 14637
rect 20416 14619 20435 14637
rect 20453 14619 20466 14637
rect 20484 14619 20494 14637
rect 19729 14613 20494 14619
rect 19729 14612 20489 14613
rect 19335 14574 19343 14592
rect 19361 14574 19369 14592
rect 19335 14553 19369 14574
rect 19335 14535 19343 14553
rect 19361 14535 19369 14553
rect 19335 14515 19369 14535
rect 19335 14497 19343 14515
rect 19361 14497 19369 14515
rect 19335 14477 19369 14497
rect 19335 14459 19343 14477
rect 19361 14459 19369 14477
rect 19335 14450 19369 14459
rect 19273 14428 19307 14434
rect 19156 14425 19307 14428
rect 18913 14392 18950 14410
rect 19156 14407 19281 14425
rect 19299 14407 19307 14425
rect 19156 14404 19307 14407
rect 19273 14398 19307 14404
rect 19343 14408 19361 14450
rect 18932 14324 18950 14392
rect 19343 14390 19392 14408
rect 18976 14324 19206 14329
rect 19374 14324 19392 14390
rect 18932 14323 19392 14324
rect 18932 14306 18988 14323
rect 18976 14305 18988 14306
rect 19006 14305 19039 14323
rect 19057 14305 19085 14323
rect 19103 14305 19131 14323
rect 19149 14305 19175 14323
rect 19193 14306 19392 14323
rect 19193 14305 19206 14306
rect 18976 14297 19206 14305
rect 17908 13931 18360 13949
rect 17353 13823 17387 13831
rect 17353 13805 17361 13823
rect 17379 13805 17387 13823
rect 17353 13785 17387 13805
rect 17353 13767 17361 13785
rect 17379 13767 17387 13785
rect 17353 13747 17387 13767
rect 17353 13729 17361 13747
rect 17379 13729 17387 13747
rect 17353 13708 17387 13729
rect 17353 13690 17361 13708
rect 17379 13690 17387 13708
rect 17353 13664 17387 13690
rect 17353 13646 17361 13664
rect 17379 13646 17387 13664
rect 17353 13626 17387 13646
rect 17353 13608 17361 13626
rect 17379 13608 17387 13626
rect 17353 13585 17387 13608
rect 17353 13567 17361 13585
rect 17379 13567 17387 13585
rect 17353 13547 17387 13567
rect 17353 13529 17361 13547
rect 17379 13529 17387 13547
rect 17353 13508 17387 13529
rect 17353 13490 17361 13508
rect 17379 13490 17387 13508
rect 17353 13467 17387 13490
rect 17353 13449 17361 13467
rect 17379 13449 17387 13467
rect 17353 13434 17387 13449
rect 17425 13823 17459 13832
rect 17908 13831 17929 13931
rect 17963 13876 17997 13885
rect 17963 13858 17971 13876
rect 17989 13858 19101 13876
rect 17963 13849 17997 13858
rect 17425 13805 17433 13823
rect 17451 13805 17459 13823
rect 17425 13785 17459 13805
rect 17425 13767 17433 13785
rect 17451 13767 17459 13785
rect 17425 13747 17459 13767
rect 17425 13729 17433 13747
rect 17451 13729 17459 13747
rect 17425 13708 17459 13729
rect 17425 13690 17433 13708
rect 17451 13690 17459 13708
rect 17425 13664 17459 13690
rect 17425 13646 17433 13664
rect 17451 13646 17459 13664
rect 17425 13626 17459 13646
rect 17425 13608 17433 13626
rect 17451 13608 17459 13626
rect 17425 13585 17459 13608
rect 17425 13567 17433 13585
rect 17451 13567 17459 13585
rect 17425 13547 17459 13567
rect 17425 13529 17433 13547
rect 17451 13529 17459 13547
rect 17425 13508 17459 13529
rect 17425 13490 17433 13508
rect 17451 13490 17459 13508
rect 17425 13467 17459 13490
rect 17425 13449 17433 13467
rect 17451 13449 17459 13467
rect 17425 13434 17459 13449
rect 17901 13823 17935 13831
rect 17901 13805 17909 13823
rect 17927 13805 17935 13823
rect 17901 13785 17935 13805
rect 17901 13767 17909 13785
rect 17927 13767 17935 13785
rect 17901 13747 17935 13767
rect 17901 13729 17909 13747
rect 17927 13729 17935 13747
rect 17901 13708 17935 13729
rect 17901 13690 17909 13708
rect 17927 13690 17935 13708
rect 17901 13664 17935 13690
rect 17901 13646 17909 13664
rect 17927 13646 17935 13664
rect 17901 13626 17935 13646
rect 17901 13608 17909 13626
rect 17927 13608 17935 13626
rect 17901 13585 17935 13608
rect 17901 13567 17909 13585
rect 17927 13567 17935 13585
rect 17901 13547 17935 13567
rect 17901 13529 17909 13547
rect 17927 13529 17935 13547
rect 17901 13508 17935 13529
rect 17901 13490 17909 13508
rect 17927 13490 17935 13508
rect 17901 13467 17935 13490
rect 17901 13449 17909 13467
rect 17927 13449 17935 13467
rect 17901 13434 17935 13449
rect 17973 13823 18007 13832
rect 17973 13805 17981 13823
rect 17999 13805 18007 13823
rect 17973 13785 18007 13805
rect 17973 13767 17981 13785
rect 17999 13767 18007 13785
rect 17973 13747 18007 13767
rect 17973 13729 17981 13747
rect 17999 13729 18007 13747
rect 17973 13708 18007 13729
rect 17973 13690 17981 13708
rect 17999 13690 18007 13708
rect 17973 13664 18007 13690
rect 17973 13646 17981 13664
rect 17999 13646 18007 13664
rect 17973 13626 18007 13646
rect 17973 13608 17981 13626
rect 17999 13608 18007 13626
rect 17973 13585 18007 13608
rect 17973 13567 17981 13585
rect 17999 13567 18007 13585
rect 17973 13547 18007 13567
rect 17973 13529 17981 13547
rect 17999 13529 18007 13547
rect 17973 13508 18007 13529
rect 17973 13490 17981 13508
rect 17999 13490 18007 13508
rect 17973 13467 18007 13490
rect 17973 13449 17981 13467
rect 17999 13449 18007 13467
rect 17973 13434 18007 13449
rect 17361 13385 17379 13434
rect 17981 13385 17999 13434
rect 17361 13367 17999 13385
rect 17637 13318 17655 13367
rect 17629 13310 17663 13318
rect 17629 13292 17637 13310
rect 17655 13292 17663 13310
rect 17629 13272 17663 13292
rect 17629 13254 17637 13272
rect 17655 13254 17663 13272
rect 17629 13234 17663 13254
rect 17629 13216 17637 13234
rect 17655 13216 17663 13234
rect 17629 13195 17663 13216
rect 17629 13177 17637 13195
rect 17655 13177 17663 13195
rect 17629 13154 17663 13177
rect 17629 13136 17637 13154
rect 17655 13136 17663 13154
rect 17629 13121 17663 13136
rect 17701 13310 17735 13319
rect 17701 13292 17709 13310
rect 17727 13292 17735 13310
rect 17701 13272 17735 13292
rect 17701 13254 17709 13272
rect 17727 13254 17735 13272
rect 17701 13234 17735 13254
rect 17701 13216 17709 13234
rect 17727 13216 17735 13234
rect 17701 13195 17735 13216
rect 17701 13177 17709 13195
rect 17727 13177 17735 13195
rect 17701 13154 17735 13177
rect 17701 13136 17709 13154
rect 17727 13136 17735 13154
rect 17701 13121 17735 13136
rect 17639 13089 17673 13098
rect 17639 13071 17647 13089
rect 17665 13071 17673 13089
rect 17639 13062 17673 13071
rect 17709 13022 17727 13121
rect 17577 13016 17807 13022
rect 17577 12998 17589 13016
rect 17607 12998 17640 13016
rect 17658 12998 17686 13016
rect 17704 12998 17732 13016
rect 17750 12998 17776 13016
rect 17794 12998 17807 13016
rect 17577 12990 17807 12998
rect 14203 12679 14292 12702
rect 14203 12661 14236 12679
rect 14253 12661 14292 12679
rect 14203 12640 14292 12661
rect 14236 12540 14254 12640
rect 19083 12540 19101 13858
rect 14236 12522 19101 12540
<< viali >>
rect 16256 16985 16273 17003
rect 22316 16134 22334 16151
rect 19669 15932 19687 15950
rect 19769 15932 19787 15950
rect 19890 15931 19908 15949
rect 19990 15931 20008 15949
rect 20147 15932 20165 15950
rect 20361 15932 20379 15950
rect 20448 15932 20466 15950
rect 17484 15575 17502 15593
rect 17584 15575 17602 15593
rect 17688 15575 17706 15593
rect 17780 15575 17798 15593
rect 17867 15575 17885 15593
rect 17110 15002 17128 15020
rect 17051 14798 17068 14815
rect 17537 15193 17554 15211
rect 17385 15077 17403 15095
rect 17617 15046 17634 15064
rect 17537 14999 17555 15017
rect 17812 15191 17830 15209
rect 17967 15137 17985 15155
rect 17813 14998 17831 15016
rect 17323 14799 17341 14816
rect 17562 14801 17580 14819
rect 17716 14888 17734 14906
rect 18028 14800 18045 14817
rect 17313 14482 17331 14500
rect 17417 14482 17435 14500
rect 17509 14482 17527 14500
rect 17601 14482 17619 14500
rect 17705 14482 17723 14500
rect 17797 14482 17815 14500
rect 17884 14482 17902 14500
rect 17966 14482 17984 14500
rect 18034 14482 18052 14500
rect 18880 15378 18898 15396
rect 18980 15378 18998 15396
rect 19084 15378 19102 15396
rect 19176 15378 19194 15396
rect 19263 15378 19281 15396
rect 18849 15048 18867 15065
rect 18279 15001 18297 15019
rect 18337 14800 18354 14817
rect 17277 14320 17295 14338
rect 17377 14320 17395 14338
rect 17481 14320 17499 14338
rect 17573 14320 17591 14338
rect 17660 14320 17678 14338
rect 17704 14320 17722 14338
rect 17804 14320 17822 14338
rect 17908 14320 17926 14338
rect 18000 14320 18018 14338
rect 18087 14320 18105 14338
rect 17371 13980 17389 13998
rect 17371 13858 17389 13876
rect 17972 13976 17990 13994
rect 19279 15046 19297 15063
rect 18851 14957 18869 14974
rect 18851 14410 18869 14427
rect 19281 14955 19299 14972
rect 19680 14972 19698 14989
rect 19945 14974 19963 14991
rect 20215 14974 20233 14991
rect 20486 14972 20504 14989
rect 20639 14970 20657 14988
rect 19745 14619 19763 14637
rect 19849 14619 19867 14637
rect 19941 14619 19959 14637
rect 20033 14619 20051 14637
rect 20137 14619 20155 14637
rect 20229 14619 20247 14637
rect 20316 14619 20334 14637
rect 20398 14619 20416 14637
rect 20466 14619 20484 14637
rect 19281 14408 19299 14425
rect 19039 14305 19057 14323
rect 19131 14305 19149 14323
rect 17971 13858 17989 13876
rect 17647 13071 17665 13089
rect 17640 12998 17658 13016
rect 17732 12998 17750 13016
rect 14236 12661 14253 12679
<< metal1 >>
rect 16687 17506 16739 17527
rect 16687 17480 16699 17506
rect 16725 17480 16739 17506
rect 16687 17456 16739 17480
rect 16671 17394 16760 17456
rect 16239 17076 16291 17097
rect 16239 17050 16251 17076
rect 16277 17050 16291 17076
rect 16239 17026 16291 17050
rect 16223 17003 16312 17026
rect 16223 16985 16256 17003
rect 16273 16985 16312 17003
rect 16223 16964 16312 16985
rect 16703 14675 16721 17394
rect 21334 16906 21405 16918
rect 21334 16880 21358 16906
rect 21384 16880 21405 16906
rect 21334 16866 21405 16880
rect 22295 16168 22357 16184
rect 22295 16156 22428 16168
rect 22295 16151 22381 16156
rect 22295 16134 22316 16151
rect 22334 16134 22381 16151
rect 22295 16130 22381 16134
rect 22407 16130 22428 16156
rect 22295 16116 22428 16130
rect 22295 16095 22357 16116
rect 20118 16062 21105 16090
rect 20118 16012 20146 16062
rect 20118 15956 20147 16012
rect 19653 15955 20368 15956
rect 19653 15950 20496 15955
rect 19653 15932 19669 15950
rect 19687 15932 19769 15950
rect 19787 15949 20147 15950
rect 19787 15932 19890 15949
rect 19653 15931 19890 15932
rect 19908 15931 19990 15949
rect 20008 15932 20147 15949
rect 20165 15932 20361 15950
rect 20379 15932 20448 15950
rect 20466 15932 20496 15950
rect 20008 15931 20496 15932
rect 19653 15925 20496 15931
rect 19874 15924 20032 15925
rect 20355 15924 20496 15925
rect 17659 15599 17688 15655
rect 17468 15593 17909 15599
rect 17468 15575 17484 15593
rect 17502 15575 17584 15593
rect 17602 15575 17688 15593
rect 17706 15575 17780 15593
rect 17798 15575 17867 15593
rect 17885 15575 17909 15593
rect 17468 15568 17909 15575
rect 19055 15402 19084 15458
rect 18864 15396 19305 15402
rect 18864 15378 18880 15396
rect 18898 15378 18980 15396
rect 18998 15378 19084 15396
rect 19102 15378 19176 15396
rect 19194 15378 19263 15396
rect 19281 15378 19305 15396
rect 18864 15371 19305 15378
rect 17527 15211 17563 15221
rect 17527 15193 17537 15211
rect 17554 15193 17563 15211
rect 17527 15184 17563 15193
rect 17797 15214 17849 15217
rect 17797 15187 17810 15214
rect 17836 15187 17849 15214
rect 17536 15156 17555 15184
rect 17797 15182 17849 15187
rect 17959 15156 17993 15161
rect 17536 15155 17993 15156
rect 17536 15137 17967 15155
rect 17985 15137 17993 15155
rect 17536 15135 17993 15137
rect 17959 15132 17993 15135
rect 17370 15100 17422 15103
rect 17370 15073 17383 15100
rect 17409 15073 17422 15100
rect 17370 15068 17422 15073
rect 17607 15064 17643 15074
rect 18841 15066 18875 15075
rect 18818 15065 18875 15066
rect 18818 15064 18849 15065
rect 17607 15046 17617 15064
rect 17634 15048 18849 15064
rect 18867 15048 18875 15065
rect 17634 15047 18875 15048
rect 17634 15046 17643 15047
rect 17607 15037 17643 15046
rect 18841 15038 18875 15047
rect 19272 15063 19305 15073
rect 19272 15046 19279 15063
rect 19297 15046 19305 15063
rect 19272 15036 19305 15046
rect 17102 15024 17136 15029
rect 17102 15017 17108 15024
rect 16982 14999 17108 15017
rect 17134 15017 17136 15024
rect 17529 15017 17564 15026
rect 17102 14998 17108 14999
rect 17134 14999 17537 15017
rect 17555 15016 17564 15017
rect 17805 15016 17839 15024
rect 18271 15023 18305 15028
rect 18271 15016 18277 15023
rect 17555 14999 17813 15016
rect 17134 14998 17136 14999
rect 17102 14993 17136 14998
rect 17529 14998 17813 14999
rect 17831 14998 18277 15016
rect 18303 15016 18305 15023
rect 18368 15016 18387 15017
rect 17529 14990 17564 14998
rect 17805 14990 17839 14998
rect 18271 14997 18277 14998
rect 18303 14998 18388 15016
rect 18303 14997 18305 14998
rect 18271 14992 18305 14997
rect 18368 14975 18387 14998
rect 19673 14989 19706 14999
rect 18843 14975 18877 14984
rect 18368 14974 18877 14975
rect 18368 14957 18851 14974
rect 18869 14973 18877 14974
rect 19273 14973 19307 14982
rect 18869 14972 19307 14973
rect 18869 14957 19281 14972
rect 18368 14956 19281 14957
rect 18843 14955 19281 14956
rect 19299 14955 19307 14972
rect 19673 14972 19680 14989
rect 19698 14972 19706 14989
rect 19673 14962 19706 14972
rect 19938 14991 19971 15001
rect 19938 14974 19945 14991
rect 19963 14974 19971 14991
rect 19938 14964 19971 14974
rect 20208 14991 20241 15001
rect 20208 14974 20215 14991
rect 20233 14974 20241 14991
rect 20208 14964 20241 14974
rect 20479 14989 20512 14999
rect 20631 14990 20665 14994
rect 20631 14989 20703 14990
rect 20479 14972 20486 14989
rect 20504 14972 20512 14989
rect 20479 14962 20512 14972
rect 20630 14988 20703 14989
rect 20630 14970 20639 14988
rect 20657 14970 20703 14988
rect 20630 14968 20703 14970
rect 20631 14965 20665 14968
rect 18843 14954 19307 14955
rect 18843 14947 18877 14954
rect 19273 14945 19307 14954
rect 17713 14906 17737 14912
rect 17678 14888 17716 14906
rect 17734 14888 17737 14906
rect 17044 14817 17076 14834
rect 17315 14817 17349 14826
rect 17044 14816 17349 14817
rect 17044 14815 17323 14816
rect 17044 14798 17051 14815
rect 17068 14799 17323 14815
rect 17341 14799 17349 14816
rect 17068 14798 17349 14799
rect 17044 14780 17076 14798
rect 17315 14789 17349 14798
rect 17555 14819 17590 14828
rect 17678 14819 17696 14888
rect 17713 14881 17737 14888
rect 17555 14801 17562 14819
rect 17580 14801 17696 14819
rect 18021 14821 18053 14826
rect 18021 14818 18072 14821
rect 18330 14818 18362 14836
rect 18021 14817 18362 14818
rect 17555 14792 17590 14801
rect 18021 14800 18028 14817
rect 18045 14800 18337 14817
rect 18354 14800 18362 14817
rect 18021 14796 18072 14800
rect 18021 14792 18053 14796
rect 18330 14782 18362 14800
rect 18330 14780 18361 14782
rect 17044 14778 17075 14780
rect 17044 14776 17063 14778
rect 16703 14657 16983 14675
rect 16965 14500 16983 14657
rect 19713 14637 20510 14643
rect 19706 14619 19745 14637
rect 19763 14619 19849 14637
rect 19867 14619 19941 14637
rect 19959 14619 20033 14637
rect 20051 14619 20137 14637
rect 20155 14619 20229 14637
rect 20247 14619 20316 14637
rect 20334 14619 20398 14637
rect 20416 14619 20466 14637
rect 20484 14619 20529 14637
rect 19713 14612 20510 14619
rect 20080 14562 20109 14612
rect 20457 14611 20510 14612
rect 17281 14500 18078 14506
rect 16965 14482 17313 14500
rect 17331 14482 17417 14500
rect 17435 14482 17509 14500
rect 17527 14482 17601 14500
rect 17619 14482 17705 14500
rect 17723 14482 17797 14500
rect 17815 14482 17884 14500
rect 17902 14482 17966 14500
rect 17984 14482 18034 14500
rect 18052 14482 18462 14500
rect 16965 13016 16983 14482
rect 17281 14475 18078 14482
rect 18025 14474 18078 14475
rect 17261 14338 18115 14344
rect 17261 14320 17277 14338
rect 17295 14320 17377 14338
rect 17395 14320 17481 14338
rect 17499 14320 17573 14338
rect 17591 14320 17660 14338
rect 17678 14320 17704 14338
rect 17722 14320 17804 14338
rect 17822 14320 17908 14338
rect 17926 14320 18000 14338
rect 18018 14320 18087 14338
rect 18105 14320 18115 14338
rect 17261 14313 18115 14320
rect 17363 14002 17397 14007
rect 17363 13976 17369 14002
rect 17395 13976 17397 14002
rect 17363 13971 17397 13976
rect 17964 13998 17998 14003
rect 17964 13972 17970 13998
rect 17996 13972 17998 13998
rect 17964 13967 17998 13972
rect 17363 13876 17397 13885
rect 17363 13858 17371 13876
rect 17389 13858 17397 13876
rect 17363 13849 17397 13858
rect 17963 13876 17997 13885
rect 17963 13858 17971 13876
rect 17989 13858 17997 13876
rect 17963 13849 17997 13858
rect 17639 13093 17673 13098
rect 17639 13067 17645 13093
rect 17671 13067 17673 13093
rect 17639 13062 17673 13067
rect 17577 13016 17807 13022
rect 18444 13016 18462 14482
rect 18843 14428 18877 14437
rect 18820 14427 18877 14428
rect 18820 14410 18851 14427
rect 18869 14410 18877 14427
rect 19273 14426 19307 14435
rect 18820 14409 18877 14410
rect 18843 14400 18877 14409
rect 19250 14425 19307 14426
rect 19250 14408 19281 14425
rect 19299 14408 19307 14425
rect 19250 14407 19307 14408
rect 19273 14398 19307 14407
rect 18976 14323 19206 14329
rect 18959 14305 19039 14323
rect 19057 14305 19131 14323
rect 19149 14305 19211 14323
rect 18976 14297 19206 14305
rect 19078 14242 19107 14297
rect 21077 14012 21105 16062
rect 21484 14036 21546 14052
rect 21484 14024 21617 14036
rect 21484 14020 21570 14024
rect 21415 14012 21570 14020
rect 21077 13998 21570 14012
rect 21596 13998 21617 14024
rect 21077 13984 21617 13998
rect 21415 13978 21546 13984
rect 21484 13963 21546 13978
rect 16965 12998 17640 13016
rect 17658 12998 17732 13016
rect 17750 12998 18462 13016
rect 17577 12990 17807 12998
rect 17679 12935 17708 12990
rect 14219 12752 14271 12773
rect 14219 12726 14231 12752
rect 14257 12726 14271 12752
rect 14219 12702 14271 12726
rect 14203 12679 14292 12702
rect 14203 12661 14236 12679
rect 14253 12661 14292 12679
rect 14203 12640 14292 12661
<< via1 >>
rect 16699 17480 16725 17506
rect 16251 17050 16277 17076
rect 21358 16880 21384 16906
rect 22381 16130 22407 16156
rect 17810 15209 17836 15214
rect 17810 15191 17812 15209
rect 17812 15191 17830 15209
rect 17830 15191 17836 15209
rect 17810 15187 17836 15191
rect 17383 15095 17409 15100
rect 17383 15077 17385 15095
rect 17385 15077 17403 15095
rect 17403 15077 17409 15095
rect 17383 15073 17409 15077
rect 17108 15020 17134 15024
rect 17108 15002 17110 15020
rect 17110 15002 17128 15020
rect 17128 15002 17134 15020
rect 17108 14998 17134 15002
rect 18277 15019 18303 15023
rect 18277 15001 18279 15019
rect 18279 15001 18297 15019
rect 18297 15001 18303 15019
rect 18277 14997 18303 15001
rect 17369 13998 17395 14002
rect 17369 13980 17371 13998
rect 17371 13980 17389 13998
rect 17389 13980 17395 13998
rect 17369 13976 17395 13980
rect 17970 13994 17996 13998
rect 17970 13976 17972 13994
rect 17972 13976 17990 13994
rect 17990 13976 17996 13994
rect 17970 13972 17996 13976
rect 17645 13089 17671 13093
rect 17645 13071 17647 13089
rect 17647 13071 17665 13089
rect 17665 13071 17671 13089
rect 17645 13067 17671 13071
rect 21570 13998 21596 14024
rect 14231 12726 14257 12752
<< metal2 >>
rect 16687 17507 16739 17527
rect 16687 17479 16698 17507
rect 16726 17479 16739 17507
rect 16687 17456 16739 17479
rect 16671 17394 16760 17456
rect 16239 17077 16291 17097
rect 16239 17049 16250 17077
rect 16278 17049 16291 17077
rect 16239 17026 16291 17049
rect 16223 16964 16312 17026
rect 21334 16907 21405 16918
rect 21334 16879 21357 16907
rect 21385 16879 21405 16907
rect 21334 16866 21405 16879
rect 21359 16649 21378 16866
rect 16948 16630 21378 16649
rect 16948 15020 16967 16630
rect 22295 16168 22357 16184
rect 22295 16157 22428 16168
rect 22295 16129 22380 16157
rect 22408 16129 22428 16157
rect 22295 16116 22428 16129
rect 22295 16095 22357 16116
rect 17797 15214 17849 15217
rect 17797 15187 17810 15214
rect 17836 15187 17849 15214
rect 17797 15182 17849 15187
rect 17370 15100 17422 15103
rect 17370 15073 17383 15100
rect 17409 15095 17422 15100
rect 17812 15095 17830 15182
rect 17409 15077 17830 15095
rect 17409 15073 17422 15077
rect 17370 15068 17422 15073
rect 17102 15024 17136 15029
rect 17102 15020 17108 15024
rect 16948 15001 17108 15020
rect 17102 14998 17108 15001
rect 17134 14998 17136 15024
rect 17102 14993 17136 14998
rect 18271 15023 18305 15028
rect 18271 14997 18277 15023
rect 18303 14997 18305 15023
rect 17109 13998 17128 14993
rect 18271 14992 18305 14997
rect 17363 14002 17397 14007
rect 17363 13998 17369 14002
rect 17109 13979 17369 13998
rect 17109 13089 17127 13979
rect 17363 13976 17369 13979
rect 17395 13976 17397 14002
rect 17363 13971 17397 13976
rect 17964 13998 17998 14003
rect 17964 13972 17970 13998
rect 17996 13994 17998 13998
rect 18278 13994 18297 14992
rect 17996 13975 18297 13994
rect 17996 13972 17998 13975
rect 17964 13967 17998 13972
rect 18278 13967 18297 13975
rect 21484 14036 21546 14052
rect 21484 14025 21617 14036
rect 21484 13997 21569 14025
rect 21597 13997 21617 14025
rect 21484 13984 21617 13997
rect 21484 13963 21546 13984
rect 17639 13093 17673 13098
rect 17639 13089 17645 13093
rect 17109 13071 17645 13089
rect 17639 13067 17645 13071
rect 17671 13067 17673 13093
rect 17639 13062 17673 13067
rect 14219 12753 14271 12773
rect 14219 12725 14230 12753
rect 14258 12725 14271 12753
rect 14219 12702 14271 12725
rect 14203 12640 14292 12702
<< via2 >>
rect 16698 17506 16726 17507
rect 16698 17480 16699 17506
rect 16699 17480 16725 17506
rect 16725 17480 16726 17506
rect 16698 17479 16726 17480
rect 16250 17076 16278 17077
rect 16250 17050 16251 17076
rect 16251 17050 16277 17076
rect 16277 17050 16278 17076
rect 16250 17049 16278 17050
rect 21357 16906 21385 16907
rect 21357 16880 21358 16906
rect 21358 16880 21384 16906
rect 21384 16880 21385 16906
rect 21357 16879 21385 16880
rect 22380 16156 22408 16157
rect 22380 16130 22381 16156
rect 22381 16130 22407 16156
rect 22407 16130 22408 16156
rect 22380 16129 22408 16130
rect 21569 14024 21597 14025
rect 21569 13998 21570 14024
rect 21570 13998 21596 14024
rect 21596 13998 21597 14024
rect 21569 13997 21597 13998
rect 14230 12752 14258 12753
rect 14230 12726 14231 12752
rect 14231 12726 14257 12752
rect 14257 12726 14258 12752
rect 14230 12725 14258 12726
<< metal3 >>
rect -37238 35494 -36178 35531
rect -36726 14450 -36689 35494
rect 16233 35485 17187 35522
rect -11091 35391 -10080 35428
rect -10486 17356 -10449 35391
rect 16695 17528 16732 35485
rect 39139 35384 40419 35421
rect 39694 27975 39731 35384
rect 30736 27938 39731 27975
rect 16687 17507 16739 17528
rect 16687 17479 16698 17507
rect 16726 17479 16739 17507
rect 16687 17456 16739 17479
rect 16671 17394 16760 17456
rect -10486 17319 16284 17356
rect 16247 17098 16284 17319
rect 16239 17077 16291 17098
rect 16239 17049 16250 17077
rect 16278 17049 16291 17077
rect 16239 17026 16291 17049
rect 16223 16964 16312 17026
rect 21334 16910 21406 16918
rect 30736 16910 30773 27938
rect 46591 24249 46628 24475
rect 21334 16907 30773 16910
rect 21334 16879 21357 16907
rect 21385 16879 30773 16907
rect 21334 16873 30773 16879
rect 41635 24212 46628 24249
rect 21334 16866 21406 16873
rect 22295 16168 22357 16184
rect 22295 16160 22429 16168
rect 41635 16160 41672 24212
rect 46591 23862 46628 24212
rect 22295 16157 41672 16160
rect 22295 16129 22380 16157
rect 22408 16129 41672 16157
rect 22295 16123 41672 16129
rect 22295 16116 22429 16123
rect 22295 16095 22357 16116
rect -36726 14413 14264 14450
rect 14227 12774 14264 14413
rect 21484 14036 21546 14052
rect 21484 14028 21618 14036
rect 21484 14025 37689 14028
rect 21484 13997 21569 14025
rect 21597 13997 37689 14025
rect 21484 13991 37689 13997
rect 21484 13984 21618 13991
rect 21484 13963 21546 13984
rect 14219 12753 14271 12774
rect 14219 12725 14230 12753
rect 14258 12725 14271 12753
rect 14219 12702 14271 12725
rect 14203 12640 14292 12702
rect 37652 5197 37689 13991
rect 46656 5197 46693 5602
rect 37652 5160 46693 5197
rect 46656 4483 46693 5160
<< labels >>
flabel locali s 17740 15180 17740 15180 0 FreeSans 300 0 0 0 Out2
port 1 nsew
flabel metal1 s 17554 15147 17554 15147 0 FreeSans 100 0 0 0 a1
port 2 nsew
flabel metal2 s 17817 15085 17817 15085 0 FreeSans 100 0 0 0 a2
port 3 nsew
flabel locali s 17440 13940 17440 13940 0 FreeSans 100 0 0 0 a3
port 4 nsew
flabel locali s 17915 13940 17915 13940 0 FreeSans 100 0 0 0 a4
port 5 nsew
flabel locali s 17643 13376 17643 13376 0 FreeSans 100 0 0 0 a5
port 6 nsew
flabel metal1 s 17614 14809 17614 14809 0 FreeSans 100 0 0 0 Out2
port 1 nsew
flabel locali s 17625 15184 17625 15184 0 FreeSans 300 0 0 0 Out1
port 7 nsew
flabel locali s 17741 14809 17741 14809 0 FreeSans 100 0 0 0 Out1
port 7 nsew
flabel locali s 19472 14982 19472 14982 0 FreeSans 300 0 0 0 tpsc_out
port 8 nsew
flabel locali s 19164 14815 19164 14815 0 FreeSans 100 0 0 0 t1
port 9 nsew
flabel locali s 18850 14697 18850 14697 0 FreeSans 100 0 0 0 t3
port 10 nsew
flabel locali s 19759 14984 19759 14984 0 FreeSans 100 0 0 0 b1
port 11 nsew
flabel locali s 20018 14976 20018 14976 0 FreeSans 100 0 0 0 b2
port 12 nsew
flabel locali s 20291 14976 20291 14976 0 FreeSans 100 0 0 0 b3
port 13 nsew
flabel locali s 19278 14685 19278 14685 0 FreeSans 100 0 0 0 t2
port 14 nsew
flabel metal3 s 22366 16143 22366 16143 0 FreeSans 300 0 0 0 io_analog[0]
port 15 nsew
flabel metal3 s 21347 16892 21347 16892 0 FreeSans 300 0 0 0 io_analog[1]
port 16 nsew
flabel metal3 s 16713 17424 16713 17424 0 FreeSans 300 0 0 0 vssa1
port 17 nsew
flabel metal3 s 21513 14003 21513 14003 0 FreeSans 300 0 0 0 vccd1
port 18 nsew
flabel metal3 s 14243 12645 14248 12646 0 FreeSans 300 0 0 0 io_analog[3]
port 19 nsew
flabel metal3 16266 16973 16266 16973 0 FreeSans 240 0 0 0 io_analog[2]
<< end >>
